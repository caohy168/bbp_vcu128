`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: htgd_thz
// Engineer: caohuiyang
// 
// Create Date: 2020/02/29 16:51:42
// Design Name: 
// Module Name: qam64-1024
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module qam(
input clk,reset,

input s_axis_input_tvalid,
output logic s_axis_input_tready,
input [7:0]s_axis_input_tdata,
input s_axis_input_tlast,

output logic m_axis_outputI_tvalid,
input  m_axis_outputI_tready,
output logic [15:0]m_axis_outputI_tdata,
output logic m_axis_outputI_tlast,
output logic m_axis_outputQ_tvalid,
input  m_axis_outputQ_tready,
output logic [15:0]m_axis_outputQ_tdata,
output logic m_axis_outputQ_tlast,

output logic m_axis_outputI_tvalid_8,
input  m_axis_outputI_tready_8,
output logic [7:0]m_axis_outputI_tdata_8,
output logic m_axis_outputI_tlast_8,
output logic m_axis_outputQ_tvalid_8,
input  m_axis_outputQ_tready_8,
output logic [7:0]m_axis_outputQ_tdata_8,
output logic m_axis_outputQ_tlast_8,

output logic m_axis_outputI_tvalid_qam256,
input  m_axis_outputI_tready_qam256,
output logic [15:0]m_axis_outputI_tdata_qam256,
output logic m_axis_outputI_tlast_qam256,
output logic m_axis_outputQ_tvalid_qam256,
input  m_axis_outputQ_tready_qam256,
output logic [15:0]m_axis_outputQ_tdata_qam256,
output logic m_axis_outputQ_tlast_qam256,

output logic m_axis_outputI_tvalid_qam1024,
input  m_axis_outputI_tready_qam1024,
output logic [15:0]m_axis_outputI_tdata_qam1024,
output logic m_axis_outputI_tlast_qam1024,
output logic m_axis_outputQ_tvalid_qam1024,
input  m_axis_outputQ_tready_qam1024,
output logic [15:0]m_axis_outputQ_tdata_qam1024,
output logic m_axis_outputQ_tlast_qam1024
);
logic m_axis_outputI_tready_qam1024,m_axis_outputQ_tready_qam1024;
assign m_axis_outputI_tready_qam1024=1;
assign m_axis_outputQ_tready_qam1024=1;

logic[15:0]tready_state; 
assign s_axis_input_tready = (tready_state==2)?0:1;
always @(posedge clk)begin
    if (reset) begin
      tready_state=0;
    end
    else begin
      case (tready_state)
         0:begin
            if (s_axis_input_tlast && s_axis_input_tvalid)
              tready_state <=1;
            else
              tready_state <=0;end
         1:begin
            if (!s_axis_input_tvalid)
            tready_state <=2;
            else
            tready_state <=1;end
         2:begin
            if(m_axis_outputI_tlast)tready_state<=0;
            else tready_state<=2;end 
      endcase
      end end
logic [15:0]axi_in_i=1;
logic [8:1]qam_input[255:1];
logic [6:1]qam64_bin[340:1];
logic [8:1]qam256_bin[255:1];
logic [10:1]qam1024_bin[204:1];

logic [1:2040]data_in=0;
logic [1:2040]data_in_1024=0;
always@(posedge clk)
    begin
        if(s_axis_input_tvalid)begin
            if(axi_in_i<255)axi_in_i<=axi_in_i+1;
            else axi_in_i<=1;
            qam_input[axi_in_i]<=s_axis_input_tdata;
            qam256_bin[axi_in_i]<=s_axis_input_tdata;
            
            data_in[8*(axi_in_i-1)+1]<=s_axis_input_tdata[7];
            data_in[8*(axi_in_i-1)+2]<=s_axis_input_tdata[6];
            data_in[8*(axi_in_i-1)+3]<=s_axis_input_tdata[5];
            data_in[8*(axi_in_i-1)+4]<=s_axis_input_tdata[4];
            data_in[8*(axi_in_i-1)+5]<=s_axis_input_tdata[3];
            data_in[8*(axi_in_i-1)+6]<=s_axis_input_tdata[2];
            data_in[8*(axi_in_i-1)+7]<=s_axis_input_tdata[1];
            data_in[8*(axi_in_i-1)+8]<=s_axis_input_tdata[0];
            
//            data_in_1024[8*(axi_in_i-1)+1]<=s_axis_input_tdata[0];
//            data_in_1024[8*(axi_in_i-1)+2]<=s_axis_input_tdata[1];
//            data_in_1024[8*(axi_in_i-1)+3]<=s_axis_input_tdata[2];
//            data_in_1024[8*(axi_in_i-1)+4]<=s_axis_input_tdata[3];
//            data_in_1024[8*(axi_in_i-1)+5]<=s_axis_input_tdata[4];
//            data_in_1024[8*(axi_in_i-1)+6]<=s_axis_input_tdata[5];
//            data_in_1024[8*(axi_in_i-1)+7]<=s_axis_input_tdata[6];
//            data_in_1024[8*(axi_in_i-1)+8]<=s_axis_input_tdata[7];

            data_in_1024[8*(axi_in_i-1)+1]<=s_axis_input_tdata[7];
            data_in_1024[8*(axi_in_i-1)+2]<=s_axis_input_tdata[6];
            data_in_1024[8*(axi_in_i-1)+3]<=s_axis_input_tdata[5];
            data_in_1024[8*(axi_in_i-1)+4]<=s_axis_input_tdata[4];
            data_in_1024[8*(axi_in_i-1)+5]<=s_axis_input_tdata[3];
            data_in_1024[8*(axi_in_i-1)+6]<=s_axis_input_tdata[2];
            data_in_1024[8*(axi_in_i-1)+7]<=s_axis_input_tdata[1];
            data_in_1024[8*(axi_in_i-1)+8]<=s_axis_input_tdata[0];
            
            end
        else axi_in_i<=1;
    end 
genvar j;
generate
    for (j = 1; j <=340; j = j + 1)begin: qam_bin_process
        always@(*)begin
            qam64_bin[j]<={data_in[6*(j-1)+1],data_in[6*(j-1)+2],data_in[6*(j-1)+3],
                         data_in[6*(j-1)+4],data_in[6*(j-1)+5],data_in[6*(j-1)+6]};
                         
//            qam1024_bin[j]<=
//                        {data_in_1024[10*(j-1)+10],data_in_1024[10*(j-1)+9],data_in_1024[10*(j-1)+8],
//                         data_in_1024[10*(j-1)+ 7],data_in_1024[10*(j-1)+6],data_in_1024[10*(j-1)+5],
//                         data_in_1024[10*(j-1)+ 4],data_in_1024[10*(j-1)+3],data_in_1024[10*(j-1)+2],
//                         data_in_1024[10*(j-1)+ 1]};

            qam1024_bin[j]<=
                        {data_in_1024[10*(j-1)+ 1],data_in_1024[10*(j-1)+2],data_in_1024[10*(j-1)+3],
                         data_in_1024[10*(j-1)+ 4],data_in_1024[10*(j-1)+5],data_in_1024[10*(j-1)+6],
                         data_in_1024[10*(j-1)+ 7],data_in_1024[10*(j-1)+8],data_in_1024[10*(j-1)+9],
                         data_in_1024[10*(j-1)+ 10]};
            end end
endgenerate
logic [6:1]gray32[1:64]={0,1,3,2,6,7,5,4,12,13,15,14,10,11,9,8,24,25,27,26,30,31,29,28,20,21,23,22,18,19,17,16,
48,49,51,50,54,55,53,52,60,61,63,62,58,59,57,56,40,41,43,42,46,47,45,44,36,37,39,38,34,35,33,32};
logic [6:1]qam64_gray_bin[340:1];
genvar i;
generate
    for (i = 1; i <=340; i = i + 1)begin: qam64_gray_bin_process
        always@(*)begin
            qam64_gray_bin[i]<=gray32[qam64_bin[i]+1];
            end end
endgenerate   
logic signed[15:0]Imodel_qam64[7:0]={-7,-5,-3,-1,1,3,5,7};
logic signed[15:0]Qmodel_qam64[7:0]={-7,-5,-3,-1,1,3,5,7};
logic signed[15:0]IEncmodel_qam64[0:63]={Imodel_qam64[7],-7,-7,-7,-7,-7,-7,-7,
                                          -5,-5,-5,-5,-5,-5,-5,-5,
                                          -1,-1,-1,-1,-1,-1,-1,-1,
                                          -3,-3,-3,-3,-3,-3,-3,-3,
                                          +7,+7,+7,+7,+7,+7,+7,+7,
                                          +5,+5,+5,+5,+5,+5,+5,+5,
                                          +1,+1,+1,+1,+1,+1,+1,+1,
                                          +3,+3,+3,+3,+3,+3,+3,+3};
logic signed[15:0]QEncmodel_qam64[0:63]={Qmodel_qam64[0],+5,+1,+3,-7,-5,-1,-3,
                                          +7,+5,+1,+3,-7,-5,-1,-3,
                                          +7,+5,+1,+3,-7,-5,-1,-3,
                                          +7,+5,+1,+3,-7,-5,-1,-3,
                                          +7,+5,+1,+3,-7,-5,-1,-3,
                                          +7,+5,+1,+3,-7,-5,-1,-3,
                                          +7,+5,+1,+3,-7,-5,-1,-3,
                                          +7,+5,+1,+3,-7,-5,-1,-3};
 
logic signed[7:0]IEncmodel_qam64_8[0:63]={-7,-7,-7,-7,-7,-7,-7,-7,
                                          -5,-5,-5,-5,-5,-5,-5,-5,
                                          -1,-1,-1,-1,-1,-1,-1,-1,
                                          -3,-3,-3,-3,-3,-3,-3,-3,
                                          +7,+7,+7,+7,+7,+7,+7,+7,
                                          +5,+5,+5,+5,+5,+5,+5,+5,
                                          +1,+1,+1,+1,+1,+1,+1,+1,
                                          +3,+3,+3,+3,+3,+3,+3,+3};
logic signed[7:0]QEncmodel_qam64_8[0:63]={+7,+5,+1,+3,-7,-5,-1,-3,
                                          +7,+5,+1,+3,-7,-5,-1,-3,
                                          +7,+5,+1,+3,-7,-5,-1,-3,
                                          +7,+5,+1,+3,-7,-5,-1,-3,
                                          +7,+5,+1,+3,-7,-5,-1,-3,
                                          +7,+5,+1,+3,-7,-5,-1,-3,
                                          +7,+5,+1,+3,-7,-5,-1,-3,
                                          +7,+5,+1,+3,-7,-5,-1,-3};
//logic signed[15:0]IQmodel[0:63][1:0]=
//{{Imodel[7],Qmodel[0]},{-7,5},{-7,1},{-7,3},{-7,-7},{-7,-5},{-7,-1},{-7,-3},
//                {-5,7},{-5,5},{-5,1},{-5,3},{-5,-7},{-5,-5},{-5,-1},{-5,-3},
//                {-1,7},{-1,5},{-1,1},{-1,3},{-1,-7},{-1,-5},{-1,-1},{-1,-3},
//                {-3,7},{-3,5},{-3,1},{-3,3},{-3,-7},{-3,-5},{-3,-1},{-3,-3},
//                {+7,7},{+7,5},{+7,1},{+7,3},{+7,-7},{+7,-5},{+7,-1},{+7,-3},
//                {+5,7},{+5,5},{+5,1},{+5,3},{+5,-7},{+5,-5},{+5,-1},{+5,-3},
//                {+1,7},{+1,5},{+1,1},{+1,3},{+1,-7},{+1,-5},{+1,-1},{+1,-3},
//                {+3,7},{+3,5},{+3,1},{+3,3},{+3,-7},{+3,-5},{+3,-1},{+3,-3}}; 
                                          
logic signed[7:0]IEncmodel_qam256[0:255]={
-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,
-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,    
 -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9,   
-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,
 -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1,    
 -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3,
 -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7,
 -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5,
 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15,
 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13,     
  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,
 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11,
  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1, 
  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,
  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,
  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5};
    
logic signed[7:0]QEncmodel_qam256[0:255]={
 15, 13,  9, 11, 1, 3, 7, 5, -15, -13, -9, -11, -1, -3, -7, -5, //-15(0-15)
 15, 13,  9, 11, 1, 3, 7, 5, -15, -13, -9,  11, -1, -3, -7, -5, //-13(16-31)
 15, 13,  9, 11, 1, 3, 7, 5, -15, -13, -9, -11, -1, -3, -7, -5, //-9(32-47)
 15, 13,  9, 11, 1, 3, 7, 5, -15, -13, -9, -11, -1, -3, -7, -5, //-11(48-63)
 15, 13,  9, 11, 1, 3, 7, 5, -15, -13, -9, -11, -1, -3, -7, -5, //-1(64-79)
 15, 13,  9, 11, 1, 3, 7, 5, -15, -13, -9, -11, -1, -3, -7, -5, //-3(80-95)
 15, 13,  9, 11, 1, 3, 7, 5, -15, -13, -9, -11, -1, -3, -7, -5, //-7(96-111)
 15, 13,  9, 11, 1, 3, 7, 5, -15, -13, -9, -11, -1, -3, -7, -5, //-5(112-127)
 15, 13,  9, 11, 1, 3, 7, 5, -15, -13, -9, -11, -1, -3, -7, -5, //15(128-143)
 15, 13,  9, 11, 1, 3, 7, 5, -15, -13, -9, -11, -1, -3, -7, -5, //13(144-159)
 15, 13,  9, 11, 1, 3, 7, 5, -15, -13, -9, -11, -1, -3, -7, -5, //9(160-175)
 15, 13,  9, 11, 1, 3, 7, 5, -15, -13, -9, -11, -1, -3, -7, -5, //11(176-191)
 15, 13,  9, 11, 1, 3, 7, 5, -15, -13, -9, -11, -1, -3, -7, -5, //1(192-207)
 15, 13,  9, 11, 1, 3, 7, 5, -15, -13, -9, -11, -1, -3, -7, -5, //3(208-223)
 15, 13,  9, 11, 1, 3, 7, 5, -15, -13, -9, -11, -1, -3, -7, -5, //7(224-239)
 15, 13,  9, 11, 1, 3, 7, 5, -15, -13, -9, -11, -1, -3, -7, -5};//5(240-255)
/*below is qam256 encode data=0:255;ans=qammod(data,256);x=real(ans);y=imag(ans)
ans =
  列 1 至 3
 -15.0000 +15.0000i -15.0000 +13.0000i -15.0000 + 9.0000i
  列 4 至 6
 -15.0000 +11.0000i -15.0000 + 1.0000i -15.0000 + 3.0000i
  列 7 至 9
 -15.0000 + 7.0000i -15.0000 + 5.0000i -15.0000 -15.0000i
  列 10 至 12
 -15.0000 -13.0000i -15.0000 - 9.0000i -15.0000 -11.0000i
  列 13 至 15
 -15.0000 - 1.0000i -15.0000 - 3.0000i -15.0000 - 7.0000i
  列 16 至 18
 -15.0000 - 5.0000i -13.0000 +15.0000i -13.0000 +13.0000i
  列 19 至 21
 -13.0000 + 9.0000i -13.0000 +11.0000i -13.0000 + 1.0000i
  列 22 至 24
 -13.0000 + 3.0000i -13.0000 + 7.0000i -13.0000 + 5.0000i
  列 25 至 27
 -13.0000 -15.0000i -13.0000 -13.0000i -13.0000 - 9.0000i
  列 28 至 30
 -13.0000 -11.0000i -13.0000 - 1.0000i -13.0000 - 3.0000i
  列 31 至 33
 -13.0000 - 7.0000i -13.0000 - 5.0000i  -9.0000 +15.0000i
  列 34 至 36
  -9.0000 +13.0000i  -9.0000 + 9.0000i  -9.0000 +11.0000i
  列 37 至 39
  -9.0000 + 1.0000i  -9.0000 + 3.0000i  -9.0000 + 7.0000i
  列 40 至 42
  -9.0000 + 5.0000i  -9.0000 -15.0000i  -9.0000 -13.0000i
  列 43 至 45
  -9.0000 - 9.0000i  -9.0000 -11.0000i  -9.0000 - 1.0000i
  列 46 至 48
  -9.0000 - 3.0000i  -9.0000 - 7.0000i  -9.0000 - 5.0000i
  列 49 至 51
 -11.0000 +15.0000i -11.0000 +13.0000i -11.0000 + 9.0000i
  列 52 至 54
 -11.0000 +11.0000i -11.0000 + 1.0000i -11.0000 + 3.0000i
  列 55 至 57
 -11.0000 + 7.0000i -11.0000 + 5.0000i -11.0000 -15.0000i
  列 58 至 60
 -11.0000 -13.0000i -11.0000 - 9.0000i -11.0000 -11.0000i
  列 61 至 63
 -11.0000 - 1.0000i -11.0000 - 3.0000i -11.0000 - 7.0000i
  列 64 至 66
 -11.0000 - 5.0000i  -1.0000 +15.0000i  -1.0000 +13.0000i
  列 67 至 69
  -1.0000 + 9.0000i  -1.0000 +11.0000i  -1.0000 + 1.0000i
  列 70 至 72
  -1.0000 + 3.0000i  -1.0000 + 7.0000i  -1.0000 + 5.0000i
  列 73 至 75
  -1.0000 -15.0000i  -1.0000 -13.0000i  -1.0000 - 9.0000i
  列 76 至 78
  -1.0000 -11.0000i  -1.0000 - 1.0000i  -1.0000 - 3.0000i
  列 79 至 81
  -1.0000 - 7.0000i  -1.0000 - 5.0000i  -3.0000 +15.0000i
  列 82 至 84
  -3.0000 +13.0000i  -3.0000 + 9.0000i  -3.0000 +11.0000i
  列 85 至 87
  -3.0000 + 1.0000i  -3.0000 + 3.0000i  -3.0000 + 7.0000i
  列 88 至 90
  -3.0000 + 5.0000i  -3.0000 -15.0000i  -3.0000 -13.0000i
  列 91 至 93
  -3.0000 - 9.0000i  -3.0000 -11.0000i  -3.0000 - 1.0000i
  列 94 至 96
  -3.0000 - 3.0000i  -3.0000 - 7.0000i  -3.0000 - 5.0000i
  列 97 至 99
  -7.0000 +15.0000i  -7.0000 +13.0000i  -7.0000 + 9.0000i
  列 100 至 102
  -7.0000 +11.0000i  -7.0000 + 1.0000i  -7.0000 + 3.0000i
  列 103 至 105
  -7.0000 + 7.0000i  -7.0000 + 5.0000i  -7.0000 -15.0000i
  列 106 至 108
  -7.0000 -13.0000i  -7.0000 - 9.0000i  -7.0000 -11.0000i
  列 109 至 111
  -7.0000 - 1.0000i  -7.0000 - 3.0000i  -7.0000 - 7.0000i
  列 112 至 114
  -7.0000 - 5.0000i  -5.0000 +15.0000i  -5.0000 +13.0000i
  列 115 至 117
  -5.0000 + 9.0000i  -5.0000 +11.0000i  -5.0000 + 1.0000i
  列 118 至 120
  -5.0000 + 3.0000i  -5.0000 + 7.0000i  -5.0000 + 5.0000i
  列 121 至 123
  -5.0000 -15.0000i  -5.0000 -13.0000i  -5.0000 - 9.0000i
  列 124 至 126
  -5.0000 -11.0000i  -5.0000 - 1.0000i  -5.0000 - 3.0000i
  列 127 至 129
  -5.0000 - 7.0000i  -5.0000 - 5.0000i  15.0000 +15.0000i
  列 130 至 132
  15.0000 +13.0000i  15.0000 + 9.0000i  15.0000 +11.0000i
  列 133 至 135
  15.0000 + 1.0000i  15.0000 + 3.0000i  15.0000 + 7.0000i
  列 136 至 138
  15.0000 + 5.0000i  15.0000 -15.0000i  15.0000 -13.0000i
  列 139 至 141
  15.0000 - 9.0000i  15.0000 -11.0000i  15.0000 - 1.0000i
  列 142 至 144
  15.0000 - 3.0000i  15.0000 - 7.0000i  15.0000 - 5.0000i
  列 145 至 147
  13.0000 +15.0000i  13.0000 +13.0000i  13.0000 + 9.0000i
  列 148 至 150
  13.0000 +11.0000i  13.0000 + 1.0000i  13.0000 + 3.0000i
  列 151 至 153
  13.0000 + 7.0000i  13.0000 + 5.0000i  13.0000 -15.0000i
  列 154 至 156
  13.0000 -13.0000i  13.0000 - 9.0000i  13.0000 -11.0000i
  列 157 至 159
  13.0000 - 1.0000i  13.0000 - 3.0000i  13.0000 - 7.0000i
  列 160 至 162
  13.0000 - 5.0000i   9.0000 +15.0000i   9.0000 +13.0000i
  列 163 至 165
   9.0000 + 9.0000i   9.0000 +11.0000i   9.0000 + 1.0000i
  列 166 至 168
   9.0000 + 3.0000i   9.0000 + 7.0000i   9.0000 + 5.0000i
  列 169 至 171
   9.0000 -15.0000i   9.0000 -13.0000i   9.0000 - 9.0000i
  列 172 至 174
   9.0000 -11.0000i   9.0000 - 1.0000i   9.0000 - 3.0000i
  列 175 至 177
   9.0000 - 7.0000i   9.0000 - 5.0000i  11.0000 +15.0000i
  列 178 至 180
  11.0000 +13.0000i  11.0000 + 9.0000i  11.0000 +11.0000i
  列 181 至 183
  11.0000 + 1.0000i  11.0000 + 3.0000i  11.0000 + 7.0000i
  列 184 至 186
  11.0000 + 5.0000i  11.0000 -15.0000i  11.0000 -13.0000i
  列 187 至 189
  11.0000 - 9.0000i  11.0000 -11.0000i  11.0000 - 1.0000i
  列 190 至 192
  11.0000 - 3.0000i  11.0000 - 7.0000i  11.0000 - 5.0000i
  列 193 至 195
   1.0000 +15.0000i   1.0000 +13.0000i   1.0000 + 9.0000i
  列 196 至 198
   1.0000 +11.0000i   1.0000 + 1.0000i   1.0000 + 3.0000i
  列 199 至 201
   1.0000 + 7.0000i   1.0000 + 5.0000i   1.0000 -15.0000i
  列 202 至 204
   1.0000 -13.0000i   1.0000 - 9.0000i   1.0000 -11.0000i
  列 205 至 207
   1.0000 - 1.0000i   1.0000 - 3.0000i   1.0000 - 7.0000i
  列 208 至 210
   1.0000 - 5.0000i   3.0000 +15.0000i   3.0000 +13.0000i
  列 211 至 213
   3.0000 + 9.0000i   3.0000 +11.0000i   3.0000 + 1.0000i
  列 214 至 216
   3.0000 + 3.0000i   3.0000 + 7.0000i   3.0000 + 5.0000i
  列 217 至 219
   3.0000 -15.0000i   3.0000 -13.0000i   3.0000 - 9.0000i
  列 220 至 222
   3.0000 -11.0000i   3.0000 - 1.0000i   3.0000 - 3.0000i
  列 223 至 225
   3.0000 - 7.0000i   3.0000 - 5.0000i   7.0000 +15.0000i
  列 226 至 228
   7.0000 +13.0000i   7.0000 + 9.0000i   7.0000 +11.0000i
  列 229 至 231
   7.0000 + 1.0000i   7.0000 + 3.0000i   7.0000 + 7.0000i
  列 232 至 234
   7.0000 + 5.0000i   7.0000 -15.0000i   7.0000 -13.0000i
  列 235 至 237
   7.0000 - 9.0000i   7.0000 -11.0000i   7.0000 - 1.0000i
  列 238 至 240
   7.0000 - 3.0000i   7.0000 - 7.0000i   7.0000 - 5.0000i
  列 241 至 243
   5.0000 +15.0000i   5.0000 +13.0000i   5.0000 + 9.0000i
  列 244 至 246
   5.0000 +11.0000i   5.0000 + 1.0000i   5.0000 + 3.0000i
  列 247 至 249
   5.0000 + 7.0000i   5.0000 + 5.0000i   5.0000 -15.0000i
  列 250 至 252
   5.0000 -13.0000i   5.0000 - 9.0000i   5.0000 -11.0000i
  列 253 至 255
   5.0000 - 1.0000i   5.0000 - 3.0000i   5.0000 - 7.0000i
  列 256
   5.0000 - 5.0000i
   */

logic signed[7:0]IEncmodel_qam1024[0:1023]={
   -31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,-31,
   -29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,-29,
   -25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,-25,
   -27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,-27,
   -17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,-17,
   -19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,-19,
   -23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,-23,
   -21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21,-21, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, -3, 
    -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, -7, 
    -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5, -5,
   -15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,-15,
   -13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13,-13, 
    -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9, -9,
   -11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11,-11, 
    31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 
    29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 
    17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 
    19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 
    23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23,
    21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21,  
     1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  1,  
     3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  3,  
     7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  7,  
     5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5,  5, 
    15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13,  
     9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9,  9, 
    11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11};
logic signed[7:0]QEncmodel_qam1024[0:1023]={
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11,
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11, 
    31, 29, 25, 27, 17, 19, 23, 21, 1, 3, 7, 5, 15, 13, 9, 11,-31,-29,-25,-27,-17,-19,-23,-21, -1, -3, -7, -5,-15,-13, -9,-11};
/*
data=0:1023
y=qammod(data,1023)
>> datai=real(y)
datai =
  列 1 至 23

   -31   -31   -31   -31   -31   -31   -31   -31   -31   -31   -31   -31   -31   -31   -31   -31   -31   -31   -31   -31   -31   -31   -31

  列 24 至 46

   -31   -31   -31   -31   -31   -31   -31   -31   -31   -29   -29   -29   -29   -29   -29   -29   -29   -29   -29   -29   -29   -29   -29

  列 47 至 69

   -29   -29   -29   -29   -29   -29   -29   -29   -29   -29   -29   -29   -29   -29   -29   -29   -29   -29   -25   -25   -25   -25   -25

  列 70 至 92

   -25   -25   -25   -25   -25   -25   -25   -25   -25   -25   -25   -25   -25   -25   -25   -25   -25   -25   -25   -25   -25   -25   -25

  列 93 至 115

   -25   -25   -25   -25   -27   -27   -27   -27   -27   -27   -27   -27   -27   -27   -27   -27   -27   -27   -27   -27   -27   -27   -27

  列 116 至 138

   -27   -27   -27   -27   -27   -27   -27   -27   -27   -27   -27   -27   -27   -17   -17   -17   -17   -17   -17   -17   -17   -17   -17

  列 139 至 161

   -17   -17   -17   -17   -17   -17   -17   -17   -17   -17   -17   -17   -17   -17   -17   -17   -17   -17   -17   -17   -17   -17   -19

  列 162 至 184

   -19   -19   -19   -19   -19   -19   -19   -19   -19   -19   -19   -19   -19   -19   -19   -19   -19   -19   -19   -19   -19   -19   -19

  列 185 至 207

   -19   -19   -19   -19   -19   -19   -19   -19   -23   -23   -23   -23   -23   -23   -23   -23   -23   -23   -23   -23   -23   -23   -23

  列 208 至 230

   -23   -23   -23   -23   -23   -23   -23   -23   -23   -23   -23   -23   -23   -23   -23   -23   -23   -21   -21   -21   -21   -21   -21

  列 231 至 253

   -21   -21   -21   -21   -21   -21   -21   -21   -21   -21   -21   -21   -21   -21   -21   -21   -21   -21   -21   -21   -21   -21   -21

  列 254 至 276

   -21   -21   -21    -1    -1    -1    -1    -1    -1    -1    -1    -1    -1    -1    -1    -1    -1    -1    -1    -1    -1    -1    -1

  列 277 至 299

    -1    -1    -1    -1    -1    -1    -1    -1    -1    -1    -1    -1    -3    -3    -3    -3    -3    -3    -3    -3    -3    -3    -3

  列 300 至 322

    -3    -3    -3    -3    -3    -3    -3    -3    -3    -3    -3    -3    -3    -3    -3    -3    -3    -3    -3    -3    -3    -7    -7

  列 323 至 345

    -7    -7    -7    -7    -7    -7    -7    -7    -7    -7    -7    -7    -7    -7    -7    -7    -7    -7    -7    -7    -7    -7    -7

  列 346 至 368

    -7    -7    -7    -7    -7    -7    -7    -5    -5    -5    -5    -5    -5    -5    -5    -5    -5    -5    -5    -5    -5    -5    -5

  列 369 至 391

    -5    -5    -5    -5    -5    -5    -5    -5    -5    -5    -5    -5    -5    -5    -5    -5   -15   -15   -15   -15   -15   -15   -15

  列 392 至 414

   -15   -15   -15   -15   -15   -15   -15   -15   -15   -15   -15   -15   -15   -15   -15   -15   -15   -15   -15   -15   -15   -15   -15

  列 415 至 437

   -15   -15   -13   -13   -13   -13   -13   -13   -13   -13   -13   -13   -13   -13   -13   -13   -13   -13   -13   -13   -13   -13   -13

  列 438 至 460

   -13   -13   -13   -13   -13   -13   -13   -13   -13   -13   -13    -9    -9    -9    -9    -9    -9    -9    -9    -9    -9    -9    -9

  列 461 至 483

    -9    -9    -9    -9    -9    -9    -9    -9    -9    -9    -9    -9    -9    -9    -9    -9    -9    -9    -9    -9   -11   -11   -11

  列 484 至 506

   -11   -11   -11   -11   -11   -11   -11   -11   -11   -11   -11   -11   -11   -11   -11   -11   -11   -11   -11   -11   -11   -11   -11

  列 507 至 529

   -11   -11   -11   -11   -11   -11    31    31    31    31    31    31    31    31    31    31    31    31    31    31    31    31    31

  列 530 至 552

    31    31    31    31    31    31    31    31    31    31    31    31    31    31    31    29    29    29    29    29    29    29    29

  列 553 至 575

    29    29    29    29    29    29    29    29    29    29    29    29    29    29    29    29    29    29    29    29    29    29    29

  列 576 至 598

    29    25    25    25    25    25    25    25    25    25    25    25    25    25    25    25    25    25    25    25    25    25    25

  列 599 至 621

    25    25    25    25    25    25    25    25    25    25    27    27    27    27    27    27    27    27    27    27    27    27    27

  列 622 至 644

    27    27    27    27    27    27    27    27    27    27    27    27    27    27    27    27    27    27    27    17    17    17    17

  列 645 至 667

    17    17    17    17    17    17    17    17    17    17    17    17    17    17    17    17    17    17    17    17    17    17    17

  列 668 至 690

    17    17    17    17    17    19    19    19    19    19    19    19    19    19    19    19    19    19    19    19    19    19    19

  列 691 至 713

    19    19    19    19    19    19    19    19    19    19    19    19    19    19    23    23    23    23    23    23    23    23    23

  列 714 至 736

    23    23    23    23    23    23    23    23    23    23    23    23    23    23    23    23    23    23    23    23    23    23    23

  列 737 至 759

    21    21    21    21    21    21    21    21    21    21    21    21    21    21    21    21    21    21    21    21    21    21    21

  列 760 至 782

    21    21    21    21    21    21    21    21    21     1     1     1     1     1     1     1     1     1     1     1     1     1     1

  列 783 至 805

     1     1     1     1     1     1     1     1     1     1     1     1     1     1     1     1     1     1     3     3     3     3     3

  列 806 至 828

     3     3     3     3     3     3     3     3     3     3     3     3     3     3     3     3     3     3     3     3     3     3     3

  列 829 至 851

     3     3     3     3     7     7     7     7     7     7     7     7     7     7     7     7     7     7     7     7     7     7     7

  列 852 至 874

     7     7     7     7     7     7     7     7     7     7     7     7     7     5     5     5     5     5     5     5     5     5     5

  列 875 至 897

     5     5     5     5     5     5     5     5     5     5     5     5     5     5     5     5     5     5     5     5     5     5    15

  列 898 至 920

    15    15    15    15    15    15    15    15    15    15    15    15    15    15    15    15    15    15    15    15    15    15    15

  列 921 至 943

    15    15    15    15    15    15    15    15    13    13    13    13    13    13    13    13    13    13    13    13    13    13    13

  列 944 至 966

    13    13    13    13    13    13    13    13    13    13    13    13    13    13    13    13    13     9     9     9     9     9     9

  列 967 至 989

     9     9     9     9     9     9     9     9     9     9     9     9     9     9     9     9     9     9     9     9     9     9     9

  列 990 至 1012

     9     9     9    11    11    11    11    11    11    11    11    11    11    11    11    11    11    11    11    11    11    11    11

  列 1013 至 1024

    11    11    11    11    11    11    11    11    11    11    11    11

>> dataq=imag(y)

dataq =

  列 1 至 23

    31    29    25    27    17    19    23    21     1     3     7     5    15    13     9    11   -31   -29   -25   -27   -17   -19   -23

  列 24 至 46

   -21    -1    -3    -7    -5   -15   -13    -9   -11    31    29    25    27    17    19    23    21     1     3     7     5    15    13

  列 47 至 69

     9    11   -31   -29   -25   -27   -17   -19   -23   -21    -1    -3    -7    -5   -15   -13    -9   -11    31    29    25    27    17

  列 70 至 92

    19    23    21     1     3     7     5    15    13     9    11   -31   -29   -25   -27   -17   -19   -23   -21    -1    -3    -7    -5

  列 93 至 115

   -15   -13    -9   -11    31    29    25    27    17    19    23    21     1     3     7     5    15    13     9    11   -31   -29   -25

  列 116 至 138

   -27   -17   -19   -23   -21    -1    -3    -7    -5   -15   -13    -9   -11    31    29    25    27    17    19    23    21     1     3

  列 139 至 161

     7     5    15    13     9    11   -31   -29   -25   -27   -17   -19   -23   -21    -1    -3    -7    -5   -15   -13    -9   -11    31

  列 162 至 184

    29    25    27    17    19    23    21     1     3     7     5    15    13     9    11   -31   -29   -25   -27   -17   -19   -23   -21

  列 185 至 207

    -1    -3    -7    -5   -15   -13    -9   -11    31    29    25    27    17    19    23    21     1     3     7     5    15    13     9

  列 208 至 230

    11   -31   -29   -25   -27   -17   -19   -23   -21    -1    -3    -7    -5   -15   -13    -9   -11    31    29    25    27    17    19

  列 231 至 253

    23    21     1     3     7     5    15    13     9    11   -31   -29   -25   -27   -17   -19   -23   -21    -1    -3    -7    -5   -15

  列 254 至 276

   -13    -9   -11    31    29    25    27    17    19    23    21     1     3     7     5    15    13     9    11   -31   -29   -25   -27

  列 277 至 299

   -17   -19   -23   -21    -1    -3    -7    -5   -15   -13    -9   -11    31    29    25    27    17    19    23    21     1     3     7

  列 300 至 322

     5    15    13     9    11   -31   -29   -25   -27   -17   -19   -23   -21    -1    -3    -7    -5   -15   -13    -9   -11    31    29

  列 323 至 345

    25    27    17    19    23    21     1     3     7     5    15    13     9    11   -31   -29   -25   -27   -17   -19   -23   -21    -1

  列 346 至 368

    -3    -7    -5   -15   -13    -9   -11    31    29    25    27    17    19    23    21     1     3     7     5    15    13     9    11

  列 369 至 391

   -31   -29   -25   -27   -17   -19   -23   -21    -1    -3    -7    -5   -15   -13    -9   -11    31    29    25    27    17    19    23

  列 392 至 414

    21     1     3     7     5    15    13     9    11   -31   -29   -25   -27   -17   -19   -23   -21    -1    -3    -7    -5   -15   -13

  列 415 至 437

    -9   -11    31    29    25    27    17    19    23    21     1     3     7     5    15    13     9    11   -31   -29   -25   -27   -17

  列 438 至 460

   -19   -23   -21    -1    -3    -7    -5   -15   -13    -9   -11    31    29    25    27    17    19    23    21     1     3     7     5

  列 461 至 483

    15    13     9    11   -31   -29   -25   -27   -17   -19   -23   -21    -1    -3    -7    -5   -15   -13    -9   -11    31    29    25

  列 484 至 506

    27    17    19    23    21     1     3     7     5    15    13     9    11   -31   -29   -25   -27   -17   -19   -23   -21    -1    -3

  列 507 至 529

    -7    -5   -15   -13    -9   -11    31    29    25    27    17    19    23    21     1     3     7     5    15    13     9    11   -31

  列 530 至 552

   -29   -25   -27   -17   -19   -23   -21    -1    -3    -7    -5   -15   -13    -9   -11    31    29    25    27    17    19    23    21

  列 553 至 575

     1     3     7     5    15    13     9    11   -31   -29   -25   -27   -17   -19   -23   -21    -1    -3    -7    -5   -15   -13    -9

  列 576 至 598

   -11    31    29    25    27    17    19    23    21     1     3     7     5    15    13     9    11   -31   -29   -25   -27   -17   -19

  列 599 至 621

   -23   -21    -1    -3    -7    -5   -15   -13    -9   -11    31    29    25    27    17    19    23    21     1     3     7     5    15

  列 622 至 644

    13     9    11   -31   -29   -25   -27   -17   -19   -23   -21    -1    -3    -7    -5   -15   -13    -9   -11    31    29    25    27

  列 645 至 667

    17    19    23    21     1     3     7     5    15    13     9    11   -31   -29   -25   -27   -17   -19   -23   -21    -1    -3    -7

  列 668 至 690

    -5   -15   -13    -9   -11    31    29    25    27    17    19    23    21     1     3     7     5    15    13     9    11   -31   -29

  列 691 至 713

   -25   -27   -17   -19   -23   -21    -1    -3    -7    -5   -15   -13    -9   -11    31    29    25    27    17    19    23    21     1

  列 714 至 736

     3     7     5    15    13     9    11   -31   -29   -25   -27   -17   -19   -23   -21    -1    -3    -7    -5   -15   -13    -9   -11

  列 737 至 759

    31    29    25    27    17    19    23    21     1     3     7     5    15    13     9    11   -31   -29   -25   -27   -17   -19   -23

  列 760 至 782

   -21    -1    -3    -7    -5   -15   -13    -9   -11    31    29    25    27    17    19    23    21     1     3     7     5    15    13

  列 783 至 805

     9    11   -31   -29   -25   -27   -17   -19   -23   -21    -1    -3    -7    -5   -15   -13    -9   -11    31    29    25    27    17

  列 806 至 828

    19    23    21     1     3     7     5    15    13     9    11   -31   -29   -25   -27   -17   -19   -23   -21    -1    -3    -7    -5

  列 829 至 851

   -15   -13    -9   -11    31    29    25    27    17    19    23    21     1     3     7     5    15    13     9    11   -31   -29   -25

  列 852 至 874

   -27   -17   -19   -23   -21    -1    -3    -7    -5   -15   -13    -9   -11    31    29    25    27    17    19    23    21     1     3

  列 875 至 897

     7     5    15    13     9    11   -31   -29   -25   -27   -17   -19   -23   -21    -1    -3    -7    -5   -15   -13    -9   -11    31

  列 898 至 920

    29    25    27    17    19    23    21     1     3     7     5    15    13     9    11   -31   -29   -25   -27   -17   -19   -23   -21

  列 921 至 943

    -1    -3    -7    -5   -15   -13    -9   -11    31    29    25    27    17    19    23    21     1     3     7     5    15    13     9

  列 944 至 966

    11   -31   -29   -25   -27   -17   -19   -23   -21    -1    -3    -7    -5   -15   -13    -9   -11    31    29    25    27    17    19

  列 967 至 989

    23    21     1     3     7     5    15    13     9    11   -31   -29   -25   -27   -17   -19   -23   -21    -1    -3    -7    -5   -15

  列 990 至 1012

   -13    -9   -11    31    29    25    27    17    19    23    21     1     3     7     5    15    13     9    11   -31   -29   -25   -27

  列 1013 至 1024

   -17   -19   -23   -21    -1    -3    -7    -5   -15   -13    -9   -11*/

logic signed[15:0]Isymbol_qam64[340:1];
logic signed[15:0]Qsymbol_qam64[340:1];
logic signed[7:0]Isymbol_qam64_8[340:1];
logic signed[7:0]Qsymbol_qam64_8[340:1];
genvar k;
generate
    for (k =1 ; k <=340; k = k + 1)begin: qam64_process
        always@(*)begin
            Isymbol_qam64[k]<=IEncmodel_qam64[qam64_gray_bin[k]];
            Qsymbol_qam64[k]<=QEncmodel_qam64[qam64_gray_bin[k]];
            
            Isymbol_qam64_8[k]<=IEncmodel_qam64_8[qam64_gray_bin[k]];
            Qsymbol_qam64_8[k]<=QEncmodel_qam64_8[qam64_gray_bin[k]];
            end end
endgenerate  

logic signed[15:0]Isymbol_qam256[255:1];
logic signed[15:0]Qsymbol_qam256[255:1];
genvar l;
generate
    for (l =1 ; l <=255; l = l + 1)begin: qam256_process
        always@(*)begin
            Isymbol_qam256[l]<=IEncmodel_qam256[qam256_bin[l]];
            Qsymbol_qam256[l]<=QEncmodel_qam256[qam256_bin[l]];
            end end
endgenerate 

logic signed[15:0]Isymbol_qam1024[204:1];
logic signed[15:0]Qsymbol_qam1024[204:1];
genvar m;
generate
    for (m =1 ; m <=204; m = m + 1)begin: qam1024_process
        always@(*)begin
            Isymbol_qam1024[m]<=IEncmodel_qam1024[qam1024_bin[m]];
            Qsymbol_qam1024[m]<=QEncmodel_qam1024[qam1024_bin[m]];
            end end
endgenerate   

logic[15:0]axi_out_i=0;  
logic[15:0]axi_out_state; 
always @(posedge clk)begin
if (reset) begin
  axi_out_state=0;
end
else begin
  case (axi_out_state)
     0: begin
        if (s_axis_input_tlast && s_axis_input_tvalid)
          axi_out_state <=1;
        else
          axi_out_state <=0;
     end
     1: begin
        if (m_axis_outputI_tready)
          axi_out_state <=2;
        else
          axi_out_state <=1;
     end
     2:begin
        if(axi_out_i<340)
            begin
                axi_out_i<=axi_out_i+1;
                axi_out_state<=2;
            end
        else begin
            axi_out_i<=0;
            axi_out_state<=0;
        end 
     end
  endcase
  end end

always@(posedge clk)
      begin
          if((axi_out_i>=1)&&(axi_out_i<=340)&&(axi_out_state==2))begin
              m_axis_outputI_tvalid<=1;
              m_axis_outputI_tdata<=Isymbol_qam64[axi_out_i];
              m_axis_outputQ_tvalid<=1;
              m_axis_outputQ_tdata<=Qsymbol_qam64[axi_out_i];
              end
          else begin
              m_axis_outputI_tvalid<=0;
              m_axis_outputI_tdata<=0;
              m_axis_outputQ_tvalid<=0;
              m_axis_outputQ_tdata<=0;
              end
          if((axi_out_i==340)&&(axi_out_state==2))m_axis_outputI_tlast<=1;
          else m_axis_outputI_tlast<=0;
          if((axi_out_i==340)&&(axi_out_state==2))m_axis_outputQ_tlast<=1;
          else m_axis_outputQ_tlast<=0;
      end
  
logic[15:0]axi_out_i_8=0;  
logic[15:0]axi_out_state_8; 
always @(posedge clk)begin
if (reset) begin
  axi_out_state_8=0;
end
else begin
  case (axi_out_state)
     0: begin
        if (s_axis_input_tlast && s_axis_input_tvalid)
          axi_out_state_8 <=1;
        else
          axi_out_state_8 <=0;
     end
     1: begin
        if (m_axis_outputI_tready_8)
          axi_out_state_8 <=2;
        else
          axi_out_state_8 <=1;
     end
     2:begin
        if(axi_out_i_8<340)
            begin
                axi_out_i_8<=axi_out_i_8+1;
                axi_out_state_8<=2;
            end
        else begin
            axi_out_i_8<=0;
            axi_out_state_8<=0;
        end 
     end
  endcase
  end end  
      
 always@(posedge clk)
      begin
          if((axi_out_i_8>=1)&&(axi_out_i_8<=340)&&(axi_out_state_8==2))begin
              m_axis_outputI_tvalid_8<=1;
              m_axis_outputI_tdata_8<=Isymbol_qam64_8[axi_out_i];
              m_axis_outputQ_tvalid_8<=1;
              m_axis_outputQ_tdata_8<=Qsymbol_qam64_8[axi_out_i];
              end
          else begin
              m_axis_outputI_tvalid_8<=0;
              m_axis_outputI_tdata_8<=0;
              m_axis_outputQ_tvalid_8<=0;
              m_axis_outputQ_tdata_8<=0;
              end
          if((axi_out_i_8==340)&&(axi_out_state_8==2))m_axis_outputI_tlast_8<=1;
          else m_axis_outputI_tlast_8<=0;
          if((axi_out_i_8==340)&&(axi_out_state_8==2))m_axis_outputQ_tlast_8<=1;
          else m_axis_outputQ_tlast_8<=0;
      end   
      
logic[15:0]axi_out_i_qam256=0;  
logic[15:0]axi_out_state_qam256; 
always @(posedge clk)begin
if (reset) begin
  axi_out_state_qam256=0;
end
else begin
  case (axi_out_state_qam256)
     0: begin
        if (s_axis_input_tlast && s_axis_input_tvalid)
          axi_out_state_qam256 <=1;
        else
          axi_out_state_qam256 <=0;
     end
     1: begin
        if (m_axis_outputI_tready_qam256)
          axi_out_state_qam256 <=2;
        else
          axi_out_state_qam256 <=1;
     end
     2:begin
        if(axi_out_i_qam256<255)
            begin
                axi_out_i_qam256<=axi_out_i_qam256+1;
                axi_out_state_qam256<=2;
            end
        else begin
            axi_out_i_qam256<=0;
            axi_out_state_qam256<=0;
        end 
     end
  endcase
  end end

always@(posedge clk)
      begin
          if((axi_out_i_qam256>=1)&&(axi_out_i_qam256<=255)&&(axi_out_state_qam256==2))begin
              m_axis_outputI_tvalid_qam256<=1;
              m_axis_outputI_tdata_qam256<=Isymbol_qam256[axi_out_i_qam256];
              m_axis_outputQ_tvalid_qam256<=1;
              m_axis_outputQ_tdata_qam256<=Qsymbol_qam256[axi_out_i_qam256];
              end
          else begin
              m_axis_outputI_tvalid_qam256<=0;
              m_axis_outputI_tdata_qam256<=0;
              m_axis_outputQ_tvalid_qam256<=0;
              m_axis_outputQ_tdata_qam256<=0;
              end
          if((axi_out_i==255)&&(axi_out_state_qam256==2))m_axis_outputI_tlast_qam256<=1;
          else m_axis_outputI_tlast_qam256<=0;
          if((axi_out_i==255)&&(axi_out_state_qam256==2))m_axis_outputQ_tlast_qam256<=1;
          else m_axis_outputQ_tlast_qam256<=0;
      end
      
logic[15:0]axi_out_i_qam1024=0;  
logic[15:0]axi_out_state_qam1024; 
always @(posedge clk)begin
if (reset) begin
  axi_out_state_qam1024=0;
end
else begin
  case (axi_out_state_qam1024)
     0: begin
        if (s_axis_input_tlast && s_axis_input_tvalid)
          axi_out_state_qam1024 <=1;
        else
          axi_out_state_qam1024 <=0;
     end
     1: begin
        if (m_axis_outputI_tready_qam1024)
          axi_out_state_qam1024 <=2;
        else
          axi_out_state_qam1024 <=1;
     end
     2:begin
        if(axi_out_i_qam256<204)
            begin
                axi_out_i_qam1024<=axi_out_i_qam1024+1;
                axi_out_state_qam1024<=2;
            end
        else begin
            axi_out_i_qam1024<=0;
            axi_out_state_qam1024<=0;
        end 
     end
  endcase
  end end

always@(posedge clk)
      begin
          if((axi_out_i_qam1024>=1)&&(axi_out_i_qam1024<=204)&&(axi_out_state_qam1024==2))begin
              m_axis_outputI_tvalid_qam1024<=1;
              m_axis_outputI_tdata_qam1024<=Isymbol_qam1024[axi_out_i_qam1024];
              m_axis_outputQ_tvalid_qam1024<=1;
              m_axis_outputQ_tdata_qam1024<=Qsymbol_qam1024[axi_out_i_qam1024];
              end
          else begin
              m_axis_outputI_tvalid_qam1024<=0;
              m_axis_outputI_tdata_qam1024<=0;
              m_axis_outputQ_tvalid_qam1024<=0;
              m_axis_outputQ_tdata_qam1024<=0;
              end
          if((axi_out_i==204)&&(axi_out_state_qam1024==2))m_axis_outputI_tlast_qam1024<=1;
          else m_axis_outputI_tlast_qam1024<=0;
          if((axi_out_i==204)&&(axi_out_state_qam1024==2))m_axis_outputQ_tlast_qam1024<=1;
          else m_axis_outputQ_tlast_qam1024<=0;
      end
       
endmodule
