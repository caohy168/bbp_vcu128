
`include "sample_tests_r.vh"
