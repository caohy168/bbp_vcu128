`include "sample_tests_t.vh"

