
`include "sample_manager.sv"
`include "csv_file_dump.sv"
`include "df_fifo_monitor.sv"
`include "df_process_monitor.sv"
`include "nodf_module_monitor.sv"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);



    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_apskdemod.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_apskdemod.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_apskdemod.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = 1'b0;
    assign module_intf_2.ap_ready = 1'b0;
    assign module_intf_2.ap_done = 1'b0;
    assign module_intf_2.ap_continue = 1'b0;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = 1'b0;
    assign module_intf_3.ap_ready = 1'b0;
    assign module_intf_3.ap_done = 1'b0;
    assign module_intf_3.ap_continue = 1'b0;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = 1'b0;
    assign module_intf_4.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_8_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_348.ap_ready;
    assign module_intf_4.ap_done = 1'b0;
    assign module_intf_4.ap_continue = 1'b0;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;
    nodf_module_intf module_intf_5(clock,reset);
    assign module_intf_5.ap_start = 1'b0;
    assign module_intf_5.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_1_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_355.ap_ready;
    assign module_intf_5.ap_done = 1'b0;
    assign module_intf_5.ap_continue = 1'b0;
    assign module_intf_5.finish = finish;
    csv_file_dump mstatus_csv_dumper_5;
    nodf_module_monitor module_monitor_5;
    nodf_module_intf module_intf_6(clock,reset);
    assign module_intf_6.ap_start = 1'b0;
    assign module_intf_6.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_4_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_363.ap_ready;
    assign module_intf_6.ap_done = 1'b0;
    assign module_intf_6.ap_continue = 1'b0;
    assign module_intf_6.finish = finish;
    csv_file_dump mstatus_csv_dumper_6;
    nodf_module_monitor module_monitor_6;
    nodf_module_intf module_intf_7(clock,reset);
    assign module_intf_7.ap_start = 1'b0;
    assign module_intf_7.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_7_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_371.ap_ready;
    assign module_intf_7.ap_done = 1'b0;
    assign module_intf_7.ap_continue = 1'b0;
    assign module_intf_7.finish = finish;
    csv_file_dump mstatus_csv_dumper_7;
    nodf_module_monitor module_monitor_7;
    nodf_module_intf module_intf_8(clock,reset);
    assign module_intf_8.ap_start = 1'b0;
    assign module_intf_8.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_12_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_378.ap_ready;
    assign module_intf_8.ap_done = 1'b0;
    assign module_intf_8.ap_continue = 1'b0;
    assign module_intf_8.finish = finish;
    csv_file_dump mstatus_csv_dumper_8;
    nodf_module_monitor module_monitor_8;
    nodf_module_intf module_intf_9(clock,reset);
    assign module_intf_9.ap_start = 1'b0;
    assign module_intf_9.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_15_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_386.ap_ready;
    assign module_intf_9.ap_done = 1'b0;
    assign module_intf_9.ap_continue = 1'b0;
    assign module_intf_9.finish = finish;
    csv_file_dump mstatus_csv_dumper_9;
    nodf_module_monitor module_monitor_9;
    nodf_module_intf module_intf_10(clock,reset);
    assign module_intf_10.ap_start = 1'b0;
    assign module_intf_10.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_18_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_394.ap_ready;
    assign module_intf_10.ap_done = 1'b0;
    assign module_intf_10.ap_continue = 1'b0;
    assign module_intf_10.finish = finish;
    csv_file_dump mstatus_csv_dumper_10;
    nodf_module_monitor module_monitor_10;
    nodf_module_intf module_intf_11(clock,reset);
    assign module_intf_11.ap_start = 1'b0;
    assign module_intf_11.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_21_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_402.ap_ready;
    assign module_intf_11.ap_done = 1'b0;
    assign module_intf_11.ap_continue = 1'b0;
    assign module_intf_11.finish = finish;
    csv_file_dump mstatus_csv_dumper_11;
    nodf_module_monitor module_monitor_11;
    nodf_module_intf module_intf_12(clock,reset);
    assign module_intf_12.ap_start = 1'b0;
    assign module_intf_12.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_24_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_410.ap_ready;
    assign module_intf_12.ap_done = 1'b0;
    assign module_intf_12.ap_continue = 1'b0;
    assign module_intf_12.finish = finish;
    csv_file_dump mstatus_csv_dumper_12;
    nodf_module_monitor module_monitor_12;
    nodf_module_intf module_intf_13(clock,reset);
    assign module_intf_13.ap_start = 1'b0;
    assign module_intf_13.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_27_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_417.ap_ready;
    assign module_intf_13.ap_done = 1'b0;
    assign module_intf_13.ap_continue = 1'b0;
    assign module_intf_13.finish = finish;
    csv_file_dump mstatus_csv_dumper_13;
    nodf_module_monitor module_monitor_13;
    nodf_module_intf module_intf_14(clock,reset);
    assign module_intf_14.ap_start = 1'b0;
    assign module_intf_14.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_30_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_425.ap_ready;
    assign module_intf_14.ap_done = 1'b0;
    assign module_intf_14.ap_continue = 1'b0;
    assign module_intf_14.finish = finish;
    csv_file_dump mstatus_csv_dumper_14;
    nodf_module_monitor module_monitor_14;
    nodf_module_intf module_intf_15(clock,reset);
    assign module_intf_15.ap_start = 1'b0;
    assign module_intf_15.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_33_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_433.ap_ready;
    assign module_intf_15.ap_done = 1'b0;
    assign module_intf_15.ap_continue = 1'b0;
    assign module_intf_15.finish = finish;
    csv_file_dump mstatus_csv_dumper_15;
    nodf_module_monitor module_monitor_15;
    nodf_module_intf module_intf_16(clock,reset);
    assign module_intf_16.ap_start = 1'b0;
    assign module_intf_16.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_36_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_441.ap_ready;
    assign module_intf_16.ap_done = 1'b0;
    assign module_intf_16.ap_continue = 1'b0;
    assign module_intf_16.finish = finish;
    csv_file_dump mstatus_csv_dumper_16;
    nodf_module_monitor module_monitor_16;
    nodf_module_intf module_intf_17(clock,reset);
    assign module_intf_17.ap_start = 1'b0;
    assign module_intf_17.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_39_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_449.ap_ready;
    assign module_intf_17.ap_done = 1'b0;
    assign module_intf_17.ap_continue = 1'b0;
    assign module_intf_17.finish = finish;
    csv_file_dump mstatus_csv_dumper_17;
    nodf_module_monitor module_monitor_17;
    nodf_module_intf module_intf_18(clock,reset);
    assign module_intf_18.ap_start = 1'b0;
    assign module_intf_18.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_42_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_456.ap_ready;
    assign module_intf_18.ap_done = 1'b0;
    assign module_intf_18.ap_continue = 1'b0;
    assign module_intf_18.finish = finish;
    csv_file_dump mstatus_csv_dumper_18;
    nodf_module_monitor module_monitor_18;
    nodf_module_intf module_intf_19(clock,reset);
    assign module_intf_19.ap_start = 1'b0;
    assign module_intf_19.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_45_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_464.ap_ready;
    assign module_intf_19.ap_done = 1'b0;
    assign module_intf_19.ap_continue = 1'b0;
    assign module_intf_19.finish = finish;
    csv_file_dump mstatus_csv_dumper_19;
    nodf_module_monitor module_monitor_19;
    nodf_module_intf module_intf_20(clock,reset);
    assign module_intf_20.ap_start = 1'b0;
    assign module_intf_20.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_48_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_472.ap_ready;
    assign module_intf_20.ap_done = 1'b0;
    assign module_intf_20.ap_continue = 1'b0;
    assign module_intf_20.finish = finish;
    csv_file_dump mstatus_csv_dumper_20;
    nodf_module_monitor module_monitor_20;
    nodf_module_intf module_intf_21(clock,reset);
    assign module_intf_21.ap_start = 1'b0;
    assign module_intf_21.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_51_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_480.ap_ready;
    assign module_intf_21.ap_done = 1'b0;
    assign module_intf_21.ap_continue = 1'b0;
    assign module_intf_21.finish = finish;
    csv_file_dump mstatus_csv_dumper_21;
    nodf_module_monitor module_monitor_21;
    nodf_module_intf module_intf_22(clock,reset);
    assign module_intf_22.ap_start = 1'b0;
    assign module_intf_22.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_54_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_488.ap_ready;
    assign module_intf_22.ap_done = 1'b0;
    assign module_intf_22.ap_continue = 1'b0;
    assign module_intf_22.finish = finish;
    csv_file_dump mstatus_csv_dumper_22;
    nodf_module_monitor module_monitor_22;
    nodf_module_intf module_intf_23(clock,reset);
    assign module_intf_23.ap_start = 1'b0;
    assign module_intf_23.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_57_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_495.ap_ready;
    assign module_intf_23.ap_done = 1'b0;
    assign module_intf_23.ap_continue = 1'b0;
    assign module_intf_23.finish = finish;
    csv_file_dump mstatus_csv_dumper_23;
    nodf_module_monitor module_monitor_23;
    nodf_module_intf module_intf_24(clock,reset);
    assign module_intf_24.ap_start = 1'b0;
    assign module_intf_24.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_60_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_503.ap_ready;
    assign module_intf_24.ap_done = 1'b0;
    assign module_intf_24.ap_continue = 1'b0;
    assign module_intf_24.finish = finish;
    csv_file_dump mstatus_csv_dumper_24;
    nodf_module_monitor module_monitor_24;
    nodf_module_intf module_intf_25(clock,reset);
    assign module_intf_25.ap_start = 1'b0;
    assign module_intf_25.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_63_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_511.ap_ready;
    assign module_intf_25.ap_done = 1'b0;
    assign module_intf_25.ap_continue = 1'b0;
    assign module_intf_25.finish = finish;
    csv_file_dump mstatus_csv_dumper_25;
    nodf_module_monitor module_monitor_25;
    nodf_module_intf module_intf_26(clock,reset);
    assign module_intf_26.ap_start = 1'b0;
    assign module_intf_26.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_66_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_519.ap_ready;
    assign module_intf_26.ap_done = 1'b0;
    assign module_intf_26.ap_continue = 1'b0;
    assign module_intf_26.finish = finish;
    csv_file_dump mstatus_csv_dumper_26;
    nodf_module_monitor module_monitor_26;
    nodf_module_intf module_intf_27(clock,reset);
    assign module_intf_27.ap_start = 1'b0;
    assign module_intf_27.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_69_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_527.ap_ready;
    assign module_intf_27.ap_done = 1'b0;
    assign module_intf_27.ap_continue = 1'b0;
    assign module_intf_27.finish = finish;
    csv_file_dump mstatus_csv_dumper_27;
    nodf_module_monitor module_monitor_27;
    nodf_module_intf module_intf_28(clock,reset);
    assign module_intf_28.ap_start = 1'b0;
    assign module_intf_28.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_72_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_534.ap_ready;
    assign module_intf_28.ap_done = 1'b0;
    assign module_intf_28.ap_continue = 1'b0;
    assign module_intf_28.finish = finish;
    csv_file_dump mstatus_csv_dumper_28;
    nodf_module_monitor module_monitor_28;
    nodf_module_intf module_intf_29(clock,reset);
    assign module_intf_29.ap_start = 1'b0;
    assign module_intf_29.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_75_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_542.ap_ready;
    assign module_intf_29.ap_done = 1'b0;
    assign module_intf_29.ap_continue = 1'b0;
    assign module_intf_29.finish = finish;
    csv_file_dump mstatus_csv_dumper_29;
    nodf_module_monitor module_monitor_29;
    nodf_module_intf module_intf_30(clock,reset);
    assign module_intf_30.ap_start = 1'b0;
    assign module_intf_30.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_78_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_550.ap_ready;
    assign module_intf_30.ap_done = 1'b0;
    assign module_intf_30.ap_continue = 1'b0;
    assign module_intf_30.finish = finish;
    csv_file_dump mstatus_csv_dumper_30;
    nodf_module_monitor module_monitor_30;
    nodf_module_intf module_intf_31(clock,reset);
    assign module_intf_31.ap_start = 1'b0;
    assign module_intf_31.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_81_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_558.ap_ready;
    assign module_intf_31.ap_done = 1'b0;
    assign module_intf_31.ap_continue = 1'b0;
    assign module_intf_31.finish = finish;
    csv_file_dump mstatus_csv_dumper_31;
    nodf_module_monitor module_monitor_31;
    nodf_module_intf module_intf_32(clock,reset);
    assign module_intf_32.ap_start = 1'b0;
    assign module_intf_32.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_84_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_566.ap_ready;
    assign module_intf_32.ap_done = 1'b0;
    assign module_intf_32.ap_continue = 1'b0;
    assign module_intf_32.finish = finish;
    csv_file_dump mstatus_csv_dumper_32;
    nodf_module_monitor module_monitor_32;
    nodf_module_intf module_intf_33(clock,reset);
    assign module_intf_33.ap_start = 1'b0;
    assign module_intf_33.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_87_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_573.ap_ready;
    assign module_intf_33.ap_done = 1'b0;
    assign module_intf_33.ap_continue = 1'b0;
    assign module_intf_33.finish = finish;
    csv_file_dump mstatus_csv_dumper_33;
    nodf_module_monitor module_monitor_33;
    nodf_module_intf module_intf_34(clock,reset);
    assign module_intf_34.ap_start = 1'b0;
    assign module_intf_34.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_90_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_581.ap_ready;
    assign module_intf_34.ap_done = 1'b0;
    assign module_intf_34.ap_continue = 1'b0;
    assign module_intf_34.finish = finish;
    csv_file_dump mstatus_csv_dumper_34;
    nodf_module_monitor module_monitor_34;
    nodf_module_intf module_intf_35(clock,reset);
    assign module_intf_35.ap_start = 1'b0;
    assign module_intf_35.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_93_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_589.ap_ready;
    assign module_intf_35.ap_done = 1'b0;
    assign module_intf_35.ap_continue = 1'b0;
    assign module_intf_35.finish = finish;
    csv_file_dump mstatus_csv_dumper_35;
    nodf_module_monitor module_monitor_35;
    nodf_module_intf module_intf_36(clock,reset);
    assign module_intf_36.ap_start = 1'b0;
    assign module_intf_36.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_96_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_597.ap_ready;
    assign module_intf_36.ap_done = 1'b0;
    assign module_intf_36.ap_continue = 1'b0;
    assign module_intf_36.finish = finish;
    csv_file_dump mstatus_csv_dumper_36;
    nodf_module_monitor module_monitor_36;
    nodf_module_intf module_intf_37(clock,reset);
    assign module_intf_37.ap_start = 1'b0;
    assign module_intf_37.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_99_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_605.ap_ready;
    assign module_intf_37.ap_done = 1'b0;
    assign module_intf_37.ap_continue = 1'b0;
    assign module_intf_37.finish = finish;
    csv_file_dump mstatus_csv_dumper_37;
    nodf_module_monitor module_monitor_37;
    nodf_module_intf module_intf_38(clock,reset);
    assign module_intf_38.ap_start = 1'b0;
    assign module_intf_38.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_102_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_612.ap_ready;
    assign module_intf_38.ap_done = 1'b0;
    assign module_intf_38.ap_continue = 1'b0;
    assign module_intf_38.finish = finish;
    csv_file_dump mstatus_csv_dumper_38;
    nodf_module_monitor module_monitor_38;
    nodf_module_intf module_intf_39(clock,reset);
    assign module_intf_39.ap_start = 1'b0;
    assign module_intf_39.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_105_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_620.ap_ready;
    assign module_intf_39.ap_done = 1'b0;
    assign module_intf_39.ap_continue = 1'b0;
    assign module_intf_39.finish = finish;
    csv_file_dump mstatus_csv_dumper_39;
    nodf_module_monitor module_monitor_39;
    nodf_module_intf module_intf_40(clock,reset);
    assign module_intf_40.ap_start = 1'b0;
    assign module_intf_40.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_108_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_628.ap_ready;
    assign module_intf_40.ap_done = 1'b0;
    assign module_intf_40.ap_continue = 1'b0;
    assign module_intf_40.finish = finish;
    csv_file_dump mstatus_csv_dumper_40;
    nodf_module_monitor module_monitor_40;
    nodf_module_intf module_intf_41(clock,reset);
    assign module_intf_41.ap_start = 1'b0;
    assign module_intf_41.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_111_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_636.ap_ready;
    assign module_intf_41.ap_done = 1'b0;
    assign module_intf_41.ap_continue = 1'b0;
    assign module_intf_41.finish = finish;
    csv_file_dump mstatus_csv_dumper_41;
    nodf_module_monitor module_monitor_41;
    nodf_module_intf module_intf_42(clock,reset);
    assign module_intf_42.ap_start = 1'b0;
    assign module_intf_42.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_114_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_644.ap_ready;
    assign module_intf_42.ap_done = 1'b0;
    assign module_intf_42.ap_continue = 1'b0;
    assign module_intf_42.finish = finish;
    csv_file_dump mstatus_csv_dumper_42;
    nodf_module_monitor module_monitor_42;
    nodf_module_intf module_intf_43(clock,reset);
    assign module_intf_43.ap_start = 1'b0;
    assign module_intf_43.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_117_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_651.ap_ready;
    assign module_intf_43.ap_done = 1'b0;
    assign module_intf_43.ap_continue = 1'b0;
    assign module_intf_43.finish = finish;
    csv_file_dump mstatus_csv_dumper_43;
    nodf_module_monitor module_monitor_43;
    nodf_module_intf module_intf_44(clock,reset);
    assign module_intf_44.ap_start = 1'b0;
    assign module_intf_44.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_119_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_659.ap_ready;
    assign module_intf_44.ap_done = 1'b0;
    assign module_intf_44.ap_continue = 1'b0;
    assign module_intf_44.finish = finish;
    csv_file_dump mstatus_csv_dumper_44;
    nodf_module_monitor module_monitor_44;
    nodf_module_intf module_intf_45(clock,reset);
    assign module_intf_45.ap_start = 1'b0;
    assign module_intf_45.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_667.ap_ready;
    assign module_intf_45.ap_done = 1'b0;
    assign module_intf_45.ap_continue = 1'b0;
    assign module_intf_45.finish = finish;
    csv_file_dump mstatus_csv_dumper_45;
    nodf_module_monitor module_monitor_45;
    nodf_module_intf module_intf_46(clock,reset);
    assign module_intf_46.ap_start = 1'b0;
    assign module_intf_46.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_s_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_674.ap_ready;
    assign module_intf_46.ap_done = 1'b0;
    assign module_intf_46.ap_continue = 1'b0;
    assign module_intf_46.finish = finish;
    csv_file_dump mstatus_csv_dumper_46;
    nodf_module_monitor module_monitor_46;
    nodf_module_intf module_intf_47(clock,reset);
    assign module_intf_47.ap_start = 1'b0;
    assign module_intf_47.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_3_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_682.ap_ready;
    assign module_intf_47.ap_done = 1'b0;
    assign module_intf_47.ap_continue = 1'b0;
    assign module_intf_47.finish = finish;
    csv_file_dump mstatus_csv_dumper_47;
    nodf_module_monitor module_monitor_47;
    nodf_module_intf module_intf_48(clock,reset);
    assign module_intf_48.ap_start = 1'b0;
    assign module_intf_48.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_6_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_690.ap_ready;
    assign module_intf_48.ap_done = 1'b0;
    assign module_intf_48.ap_continue = 1'b0;
    assign module_intf_48.finish = finish;
    csv_file_dump mstatus_csv_dumper_48;
    nodf_module_monitor module_monitor_48;
    nodf_module_intf module_intf_49(clock,reset);
    assign module_intf_49.ap_start = 1'b0;
    assign module_intf_49.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_11_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_697.ap_ready;
    assign module_intf_49.ap_done = 1'b0;
    assign module_intf_49.ap_continue = 1'b0;
    assign module_intf_49.finish = finish;
    csv_file_dump mstatus_csv_dumper_49;
    nodf_module_monitor module_monitor_49;
    nodf_module_intf module_intf_50(clock,reset);
    assign module_intf_50.ap_start = 1'b0;
    assign module_intf_50.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_14_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_705.ap_ready;
    assign module_intf_50.ap_done = 1'b0;
    assign module_intf_50.ap_continue = 1'b0;
    assign module_intf_50.finish = finish;
    csv_file_dump mstatus_csv_dumper_50;
    nodf_module_monitor module_monitor_50;
    nodf_module_intf module_intf_51(clock,reset);
    assign module_intf_51.ap_start = 1'b0;
    assign module_intf_51.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_17_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_713.ap_ready;
    assign module_intf_51.ap_done = 1'b0;
    assign module_intf_51.ap_continue = 1'b0;
    assign module_intf_51.finish = finish;
    csv_file_dump mstatus_csv_dumper_51;
    nodf_module_monitor module_monitor_51;
    nodf_module_intf module_intf_52(clock,reset);
    assign module_intf_52.ap_start = 1'b0;
    assign module_intf_52.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_20_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_721.ap_ready;
    assign module_intf_52.ap_done = 1'b0;
    assign module_intf_52.ap_continue = 1'b0;
    assign module_intf_52.finish = finish;
    csv_file_dump mstatus_csv_dumper_52;
    nodf_module_monitor module_monitor_52;
    nodf_module_intf module_intf_53(clock,reset);
    assign module_intf_53.ap_start = 1'b0;
    assign module_intf_53.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_23_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_729.ap_ready;
    assign module_intf_53.ap_done = 1'b0;
    assign module_intf_53.ap_continue = 1'b0;
    assign module_intf_53.finish = finish;
    csv_file_dump mstatus_csv_dumper_53;
    nodf_module_monitor module_monitor_53;
    nodf_module_intf module_intf_54(clock,reset);
    assign module_intf_54.ap_start = 1'b0;
    assign module_intf_54.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_26_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_736.ap_ready;
    assign module_intf_54.ap_done = 1'b0;
    assign module_intf_54.ap_continue = 1'b0;
    assign module_intf_54.finish = finish;
    csv_file_dump mstatus_csv_dumper_54;
    nodf_module_monitor module_monitor_54;
    nodf_module_intf module_intf_55(clock,reset);
    assign module_intf_55.ap_start = 1'b0;
    assign module_intf_55.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_29_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_744.ap_ready;
    assign module_intf_55.ap_done = 1'b0;
    assign module_intf_55.ap_continue = 1'b0;
    assign module_intf_55.finish = finish;
    csv_file_dump mstatus_csv_dumper_55;
    nodf_module_monitor module_monitor_55;
    nodf_module_intf module_intf_56(clock,reset);
    assign module_intf_56.ap_start = 1'b0;
    assign module_intf_56.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_32_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_752.ap_ready;
    assign module_intf_56.ap_done = 1'b0;
    assign module_intf_56.ap_continue = 1'b0;
    assign module_intf_56.finish = finish;
    csv_file_dump mstatus_csv_dumper_56;
    nodf_module_monitor module_monitor_56;
    nodf_module_intf module_intf_57(clock,reset);
    assign module_intf_57.ap_start = 1'b0;
    assign module_intf_57.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_35_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_760.ap_ready;
    assign module_intf_57.ap_done = 1'b0;
    assign module_intf_57.ap_continue = 1'b0;
    assign module_intf_57.finish = finish;
    csv_file_dump mstatus_csv_dumper_57;
    nodf_module_monitor module_monitor_57;
    nodf_module_intf module_intf_58(clock,reset);
    assign module_intf_58.ap_start = 1'b0;
    assign module_intf_58.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_38_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_768.ap_ready;
    assign module_intf_58.ap_done = 1'b0;
    assign module_intf_58.ap_continue = 1'b0;
    assign module_intf_58.finish = finish;
    csv_file_dump mstatus_csv_dumper_58;
    nodf_module_monitor module_monitor_58;
    nodf_module_intf module_intf_59(clock,reset);
    assign module_intf_59.ap_start = 1'b0;
    assign module_intf_59.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_41_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_775.ap_ready;
    assign module_intf_59.ap_done = 1'b0;
    assign module_intf_59.ap_continue = 1'b0;
    assign module_intf_59.finish = finish;
    csv_file_dump mstatus_csv_dumper_59;
    nodf_module_monitor module_monitor_59;
    nodf_module_intf module_intf_60(clock,reset);
    assign module_intf_60.ap_start = 1'b0;
    assign module_intf_60.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_44_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_783.ap_ready;
    assign module_intf_60.ap_done = 1'b0;
    assign module_intf_60.ap_continue = 1'b0;
    assign module_intf_60.finish = finish;
    csv_file_dump mstatus_csv_dumper_60;
    nodf_module_monitor module_monitor_60;
    nodf_module_intf module_intf_61(clock,reset);
    assign module_intf_61.ap_start = 1'b0;
    assign module_intf_61.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_47_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_791.ap_ready;
    assign module_intf_61.ap_done = 1'b0;
    assign module_intf_61.ap_continue = 1'b0;
    assign module_intf_61.finish = finish;
    csv_file_dump mstatus_csv_dumper_61;
    nodf_module_monitor module_monitor_61;
    nodf_module_intf module_intf_62(clock,reset);
    assign module_intf_62.ap_start = 1'b0;
    assign module_intf_62.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_50_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_799.ap_ready;
    assign module_intf_62.ap_done = 1'b0;
    assign module_intf_62.ap_continue = 1'b0;
    assign module_intf_62.finish = finish;
    csv_file_dump mstatus_csv_dumper_62;
    nodf_module_monitor module_monitor_62;
    nodf_module_intf module_intf_63(clock,reset);
    assign module_intf_63.ap_start = 1'b0;
    assign module_intf_63.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_53_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_807.ap_ready;
    assign module_intf_63.ap_done = 1'b0;
    assign module_intf_63.ap_continue = 1'b0;
    assign module_intf_63.finish = finish;
    csv_file_dump mstatus_csv_dumper_63;
    nodf_module_monitor module_monitor_63;
    nodf_module_intf module_intf_64(clock,reset);
    assign module_intf_64.ap_start = 1'b0;
    assign module_intf_64.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_56_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_814.ap_ready;
    assign module_intf_64.ap_done = 1'b0;
    assign module_intf_64.ap_continue = 1'b0;
    assign module_intf_64.finish = finish;
    csv_file_dump mstatus_csv_dumper_64;
    nodf_module_monitor module_monitor_64;
    nodf_module_intf module_intf_65(clock,reset);
    assign module_intf_65.ap_start = 1'b0;
    assign module_intf_65.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_59_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_822.ap_ready;
    assign module_intf_65.ap_done = 1'b0;
    assign module_intf_65.ap_continue = 1'b0;
    assign module_intf_65.finish = finish;
    csv_file_dump mstatus_csv_dumper_65;
    nodf_module_monitor module_monitor_65;
    nodf_module_intf module_intf_66(clock,reset);
    assign module_intf_66.ap_start = 1'b0;
    assign module_intf_66.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_62_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_830.ap_ready;
    assign module_intf_66.ap_done = 1'b0;
    assign module_intf_66.ap_continue = 1'b0;
    assign module_intf_66.finish = finish;
    csv_file_dump mstatus_csv_dumper_66;
    nodf_module_monitor module_monitor_66;
    nodf_module_intf module_intf_67(clock,reset);
    assign module_intf_67.ap_start = 1'b0;
    assign module_intf_67.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_65_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_838.ap_ready;
    assign module_intf_67.ap_done = 1'b0;
    assign module_intf_67.ap_continue = 1'b0;
    assign module_intf_67.finish = finish;
    csv_file_dump mstatus_csv_dumper_67;
    nodf_module_monitor module_monitor_67;
    nodf_module_intf module_intf_68(clock,reset);
    assign module_intf_68.ap_start = 1'b0;
    assign module_intf_68.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_68_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_846.ap_ready;
    assign module_intf_68.ap_done = 1'b0;
    assign module_intf_68.ap_continue = 1'b0;
    assign module_intf_68.finish = finish;
    csv_file_dump mstatus_csv_dumper_68;
    nodf_module_monitor module_monitor_68;
    nodf_module_intf module_intf_69(clock,reset);
    assign module_intf_69.ap_start = 1'b0;
    assign module_intf_69.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_71_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_853.ap_ready;
    assign module_intf_69.ap_done = 1'b0;
    assign module_intf_69.ap_continue = 1'b0;
    assign module_intf_69.finish = finish;
    csv_file_dump mstatus_csv_dumper_69;
    nodf_module_monitor module_monitor_69;
    nodf_module_intf module_intf_70(clock,reset);
    assign module_intf_70.ap_start = 1'b0;
    assign module_intf_70.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_74_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_861.ap_ready;
    assign module_intf_70.ap_done = 1'b0;
    assign module_intf_70.ap_continue = 1'b0;
    assign module_intf_70.finish = finish;
    csv_file_dump mstatus_csv_dumper_70;
    nodf_module_monitor module_monitor_70;
    nodf_module_intf module_intf_71(clock,reset);
    assign module_intf_71.ap_start = 1'b0;
    assign module_intf_71.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_77_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_869.ap_ready;
    assign module_intf_71.ap_done = 1'b0;
    assign module_intf_71.ap_continue = 1'b0;
    assign module_intf_71.finish = finish;
    csv_file_dump mstatus_csv_dumper_71;
    nodf_module_monitor module_monitor_71;
    nodf_module_intf module_intf_72(clock,reset);
    assign module_intf_72.ap_start = 1'b0;
    assign module_intf_72.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_80_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_877.ap_ready;
    assign module_intf_72.ap_done = 1'b0;
    assign module_intf_72.ap_continue = 1'b0;
    assign module_intf_72.finish = finish;
    csv_file_dump mstatus_csv_dumper_72;
    nodf_module_monitor module_monitor_72;
    nodf_module_intf module_intf_73(clock,reset);
    assign module_intf_73.ap_start = 1'b0;
    assign module_intf_73.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_83_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_885.ap_ready;
    assign module_intf_73.ap_done = 1'b0;
    assign module_intf_73.ap_continue = 1'b0;
    assign module_intf_73.finish = finish;
    csv_file_dump mstatus_csv_dumper_73;
    nodf_module_monitor module_monitor_73;
    nodf_module_intf module_intf_74(clock,reset);
    assign module_intf_74.ap_start = 1'b0;
    assign module_intf_74.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_86_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_892.ap_ready;
    assign module_intf_74.ap_done = 1'b0;
    assign module_intf_74.ap_continue = 1'b0;
    assign module_intf_74.finish = finish;
    csv_file_dump mstatus_csv_dumper_74;
    nodf_module_monitor module_monitor_74;
    nodf_module_intf module_intf_75(clock,reset);
    assign module_intf_75.ap_start = 1'b0;
    assign module_intf_75.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_89_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_900.ap_ready;
    assign module_intf_75.ap_done = 1'b0;
    assign module_intf_75.ap_continue = 1'b0;
    assign module_intf_75.finish = finish;
    csv_file_dump mstatus_csv_dumper_75;
    nodf_module_monitor module_monitor_75;
    nodf_module_intf module_intf_76(clock,reset);
    assign module_intf_76.ap_start = 1'b0;
    assign module_intf_76.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_92_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_908.ap_ready;
    assign module_intf_76.ap_done = 1'b0;
    assign module_intf_76.ap_continue = 1'b0;
    assign module_intf_76.finish = finish;
    csv_file_dump mstatus_csv_dumper_76;
    nodf_module_monitor module_monitor_76;
    nodf_module_intf module_intf_77(clock,reset);
    assign module_intf_77.ap_start = 1'b0;
    assign module_intf_77.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_95_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_916.ap_ready;
    assign module_intf_77.ap_done = 1'b0;
    assign module_intf_77.ap_continue = 1'b0;
    assign module_intf_77.finish = finish;
    csv_file_dump mstatus_csv_dumper_77;
    nodf_module_monitor module_monitor_77;
    nodf_module_intf module_intf_78(clock,reset);
    assign module_intf_78.ap_start = 1'b0;
    assign module_intf_78.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_98_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_924.ap_ready;
    assign module_intf_78.ap_done = 1'b0;
    assign module_intf_78.ap_continue = 1'b0;
    assign module_intf_78.finish = finish;
    csv_file_dump mstatus_csv_dumper_78;
    nodf_module_monitor module_monitor_78;
    nodf_module_intf module_intf_79(clock,reset);
    assign module_intf_79.ap_start = 1'b0;
    assign module_intf_79.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_101_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_931.ap_ready;
    assign module_intf_79.ap_done = 1'b0;
    assign module_intf_79.ap_continue = 1'b0;
    assign module_intf_79.finish = finish;
    csv_file_dump mstatus_csv_dumper_79;
    nodf_module_monitor module_monitor_79;
    nodf_module_intf module_intf_80(clock,reset);
    assign module_intf_80.ap_start = 1'b0;
    assign module_intf_80.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_104_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_939.ap_ready;
    assign module_intf_80.ap_done = 1'b0;
    assign module_intf_80.ap_continue = 1'b0;
    assign module_intf_80.finish = finish;
    csv_file_dump mstatus_csv_dumper_80;
    nodf_module_monitor module_monitor_80;
    nodf_module_intf module_intf_81(clock,reset);
    assign module_intf_81.ap_start = 1'b0;
    assign module_intf_81.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_107_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_947.ap_ready;
    assign module_intf_81.ap_done = 1'b0;
    assign module_intf_81.ap_continue = 1'b0;
    assign module_intf_81.finish = finish;
    csv_file_dump mstatus_csv_dumper_81;
    nodf_module_monitor module_monitor_81;
    nodf_module_intf module_intf_82(clock,reset);
    assign module_intf_82.ap_start = 1'b0;
    assign module_intf_82.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_110_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_955.ap_ready;
    assign module_intf_82.ap_done = 1'b0;
    assign module_intf_82.ap_continue = 1'b0;
    assign module_intf_82.finish = finish;
    csv_file_dump mstatus_csv_dumper_82;
    nodf_module_monitor module_monitor_82;
    nodf_module_intf module_intf_83(clock,reset);
    assign module_intf_83.ap_start = 1'b0;
    assign module_intf_83.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_113_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_963.ap_ready;
    assign module_intf_83.ap_done = 1'b0;
    assign module_intf_83.ap_continue = 1'b0;
    assign module_intf_83.finish = finish;
    csv_file_dump mstatus_csv_dumper_83;
    nodf_module_monitor module_monitor_83;
    nodf_module_intf module_intf_84(clock,reset);
    assign module_intf_84.ap_start = 1'b0;
    assign module_intf_84.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_116_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_970.ap_ready;
    assign module_intf_84.ap_done = 1'b0;
    assign module_intf_84.ap_continue = 1'b0;
    assign module_intf_84.finish = finish;
    csv_file_dump mstatus_csv_dumper_84;
    nodf_module_monitor module_monitor_84;
    nodf_module_intf module_intf_85(clock,reset);
    assign module_intf_85.ap_start = 1'b0;
    assign module_intf_85.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_9_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_978.ap_ready;
    assign module_intf_85.ap_done = 1'b0;
    assign module_intf_85.ap_continue = 1'b0;
    assign module_intf_85.finish = finish;
    csv_file_dump mstatus_csv_dumper_85;
    nodf_module_monitor module_monitor_85;
    nodf_module_intf module_intf_86(clock,reset);
    assign module_intf_86.ap_start = 1'b0;
    assign module_intf_86.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_2_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_987.ap_ready;
    assign module_intf_86.ap_done = 1'b0;
    assign module_intf_86.ap_continue = 1'b0;
    assign module_intf_86.finish = finish;
    csv_file_dump mstatus_csv_dumper_86;
    nodf_module_monitor module_monitor_86;
    nodf_module_intf module_intf_87(clock,reset);
    assign module_intf_87.ap_start = 1'b0;
    assign module_intf_87.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_5_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_996.ap_ready;
    assign module_intf_87.ap_done = 1'b0;
    assign module_intf_87.ap_continue = 1'b0;
    assign module_intf_87.finish = finish;
    csv_file_dump mstatus_csv_dumper_87;
    nodf_module_monitor module_monitor_87;
    nodf_module_intf module_intf_88(clock,reset);
    assign module_intf_88.ap_start = 1'b0;
    assign module_intf_88.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_10_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1005.ap_ready;
    assign module_intf_88.ap_done = 1'b0;
    assign module_intf_88.ap_continue = 1'b0;
    assign module_intf_88.finish = finish;
    csv_file_dump mstatus_csv_dumper_88;
    nodf_module_monitor module_monitor_88;
    nodf_module_intf module_intf_89(clock,reset);
    assign module_intf_89.ap_start = 1'b0;
    assign module_intf_89.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_13_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1014.ap_ready;
    assign module_intf_89.ap_done = 1'b0;
    assign module_intf_89.ap_continue = 1'b0;
    assign module_intf_89.finish = finish;
    csv_file_dump mstatus_csv_dumper_89;
    nodf_module_monitor module_monitor_89;
    nodf_module_intf module_intf_90(clock,reset);
    assign module_intf_90.ap_start = 1'b0;
    assign module_intf_90.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_16_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1023.ap_ready;
    assign module_intf_90.ap_done = 1'b0;
    assign module_intf_90.ap_continue = 1'b0;
    assign module_intf_90.finish = finish;
    csv_file_dump mstatus_csv_dumper_90;
    nodf_module_monitor module_monitor_90;
    nodf_module_intf module_intf_91(clock,reset);
    assign module_intf_91.ap_start = 1'b0;
    assign module_intf_91.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_19_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1032.ap_ready;
    assign module_intf_91.ap_done = 1'b0;
    assign module_intf_91.ap_continue = 1'b0;
    assign module_intf_91.finish = finish;
    csv_file_dump mstatus_csv_dumper_91;
    nodf_module_monitor module_monitor_91;
    nodf_module_intf module_intf_92(clock,reset);
    assign module_intf_92.ap_start = 1'b0;
    assign module_intf_92.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_22_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1040.ap_ready;
    assign module_intf_92.ap_done = 1'b0;
    assign module_intf_92.ap_continue = 1'b0;
    assign module_intf_92.finish = finish;
    csv_file_dump mstatus_csv_dumper_92;
    nodf_module_monitor module_monitor_92;
    nodf_module_intf module_intf_93(clock,reset);
    assign module_intf_93.ap_start = 1'b0;
    assign module_intf_93.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_25_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1049.ap_ready;
    assign module_intf_93.ap_done = 1'b0;
    assign module_intf_93.ap_continue = 1'b0;
    assign module_intf_93.finish = finish;
    csv_file_dump mstatus_csv_dumper_93;
    nodf_module_monitor module_monitor_93;
    nodf_module_intf module_intf_94(clock,reset);
    assign module_intf_94.ap_start = 1'b0;
    assign module_intf_94.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_28_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1058.ap_ready;
    assign module_intf_94.ap_done = 1'b0;
    assign module_intf_94.ap_continue = 1'b0;
    assign module_intf_94.finish = finish;
    csv_file_dump mstatus_csv_dumper_94;
    nodf_module_monitor module_monitor_94;
    nodf_module_intf module_intf_95(clock,reset);
    assign module_intf_95.ap_start = 1'b0;
    assign module_intf_95.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_31_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1067.ap_ready;
    assign module_intf_95.ap_done = 1'b0;
    assign module_intf_95.ap_continue = 1'b0;
    assign module_intf_95.finish = finish;
    csv_file_dump mstatus_csv_dumper_95;
    nodf_module_monitor module_monitor_95;
    nodf_module_intf module_intf_96(clock,reset);
    assign module_intf_96.ap_start = 1'b0;
    assign module_intf_96.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_34_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1076.ap_ready;
    assign module_intf_96.ap_done = 1'b0;
    assign module_intf_96.ap_continue = 1'b0;
    assign module_intf_96.finish = finish;
    csv_file_dump mstatus_csv_dumper_96;
    nodf_module_monitor module_monitor_96;
    nodf_module_intf module_intf_97(clock,reset);
    assign module_intf_97.ap_start = 1'b0;
    assign module_intf_97.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_37_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1085.ap_ready;
    assign module_intf_97.ap_done = 1'b0;
    assign module_intf_97.ap_continue = 1'b0;
    assign module_intf_97.finish = finish;
    csv_file_dump mstatus_csv_dumper_97;
    nodf_module_monitor module_monitor_97;
    nodf_module_intf module_intf_98(clock,reset);
    assign module_intf_98.ap_start = 1'b0;
    assign module_intf_98.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_40_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1093.ap_ready;
    assign module_intf_98.ap_done = 1'b0;
    assign module_intf_98.ap_continue = 1'b0;
    assign module_intf_98.finish = finish;
    csv_file_dump mstatus_csv_dumper_98;
    nodf_module_monitor module_monitor_98;
    nodf_module_intf module_intf_99(clock,reset);
    assign module_intf_99.ap_start = 1'b0;
    assign module_intf_99.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_43_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1102.ap_ready;
    assign module_intf_99.ap_done = 1'b0;
    assign module_intf_99.ap_continue = 1'b0;
    assign module_intf_99.finish = finish;
    csv_file_dump mstatus_csv_dumper_99;
    nodf_module_monitor module_monitor_99;
    nodf_module_intf module_intf_100(clock,reset);
    assign module_intf_100.ap_start = 1'b0;
    assign module_intf_100.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_46_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1111.ap_ready;
    assign module_intf_100.ap_done = 1'b0;
    assign module_intf_100.ap_continue = 1'b0;
    assign module_intf_100.finish = finish;
    csv_file_dump mstatus_csv_dumper_100;
    nodf_module_monitor module_monitor_100;
    nodf_module_intf module_intf_101(clock,reset);
    assign module_intf_101.ap_start = 1'b0;
    assign module_intf_101.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_49_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1120.ap_ready;
    assign module_intf_101.ap_done = 1'b0;
    assign module_intf_101.ap_continue = 1'b0;
    assign module_intf_101.finish = finish;
    csv_file_dump mstatus_csv_dumper_101;
    nodf_module_monitor module_monitor_101;
    nodf_module_intf module_intf_102(clock,reset);
    assign module_intf_102.ap_start = 1'b0;
    assign module_intf_102.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_52_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1129.ap_ready;
    assign module_intf_102.ap_done = 1'b0;
    assign module_intf_102.ap_continue = 1'b0;
    assign module_intf_102.finish = finish;
    csv_file_dump mstatus_csv_dumper_102;
    nodf_module_monitor module_monitor_102;
    nodf_module_intf module_intf_103(clock,reset);
    assign module_intf_103.ap_start = 1'b0;
    assign module_intf_103.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_55_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1138.ap_ready;
    assign module_intf_103.ap_done = 1'b0;
    assign module_intf_103.ap_continue = 1'b0;
    assign module_intf_103.finish = finish;
    csv_file_dump mstatus_csv_dumper_103;
    nodf_module_monitor module_monitor_103;
    nodf_module_intf module_intf_104(clock,reset);
    assign module_intf_104.ap_start = 1'b0;
    assign module_intf_104.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_58_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1146.ap_ready;
    assign module_intf_104.ap_done = 1'b0;
    assign module_intf_104.ap_continue = 1'b0;
    assign module_intf_104.finish = finish;
    csv_file_dump mstatus_csv_dumper_104;
    nodf_module_monitor module_monitor_104;
    nodf_module_intf module_intf_105(clock,reset);
    assign module_intf_105.ap_start = 1'b0;
    assign module_intf_105.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_61_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1155.ap_ready;
    assign module_intf_105.ap_done = 1'b0;
    assign module_intf_105.ap_continue = 1'b0;
    assign module_intf_105.finish = finish;
    csv_file_dump mstatus_csv_dumper_105;
    nodf_module_monitor module_monitor_105;
    nodf_module_intf module_intf_106(clock,reset);
    assign module_intf_106.ap_start = 1'b0;
    assign module_intf_106.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_64_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1164.ap_ready;
    assign module_intf_106.ap_done = 1'b0;
    assign module_intf_106.ap_continue = 1'b0;
    assign module_intf_106.finish = finish;
    csv_file_dump mstatus_csv_dumper_106;
    nodf_module_monitor module_monitor_106;
    nodf_module_intf module_intf_107(clock,reset);
    assign module_intf_107.ap_start = 1'b0;
    assign module_intf_107.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_67_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1173.ap_ready;
    assign module_intf_107.ap_done = 1'b0;
    assign module_intf_107.ap_continue = 1'b0;
    assign module_intf_107.finish = finish;
    csv_file_dump mstatus_csv_dumper_107;
    nodf_module_monitor module_monitor_107;
    nodf_module_intf module_intf_108(clock,reset);
    assign module_intf_108.ap_start = 1'b0;
    assign module_intf_108.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_70_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1182.ap_ready;
    assign module_intf_108.ap_done = 1'b0;
    assign module_intf_108.ap_continue = 1'b0;
    assign module_intf_108.finish = finish;
    csv_file_dump mstatus_csv_dumper_108;
    nodf_module_monitor module_monitor_108;
    nodf_module_intf module_intf_109(clock,reset);
    assign module_intf_109.ap_start = 1'b0;
    assign module_intf_109.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_73_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1190.ap_ready;
    assign module_intf_109.ap_done = 1'b0;
    assign module_intf_109.ap_continue = 1'b0;
    assign module_intf_109.finish = finish;
    csv_file_dump mstatus_csv_dumper_109;
    nodf_module_monitor module_monitor_109;
    nodf_module_intf module_intf_110(clock,reset);
    assign module_intf_110.ap_start = 1'b0;
    assign module_intf_110.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_76_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1199.ap_ready;
    assign module_intf_110.ap_done = 1'b0;
    assign module_intf_110.ap_continue = 1'b0;
    assign module_intf_110.finish = finish;
    csv_file_dump mstatus_csv_dumper_110;
    nodf_module_monitor module_monitor_110;
    nodf_module_intf module_intf_111(clock,reset);
    assign module_intf_111.ap_start = 1'b0;
    assign module_intf_111.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_79_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1208.ap_ready;
    assign module_intf_111.ap_done = 1'b0;
    assign module_intf_111.ap_continue = 1'b0;
    assign module_intf_111.finish = finish;
    csv_file_dump mstatus_csv_dumper_111;
    nodf_module_monitor module_monitor_111;
    nodf_module_intf module_intf_112(clock,reset);
    assign module_intf_112.ap_start = 1'b0;
    assign module_intf_112.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_82_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1217.ap_ready;
    assign module_intf_112.ap_done = 1'b0;
    assign module_intf_112.ap_continue = 1'b0;
    assign module_intf_112.finish = finish;
    csv_file_dump mstatus_csv_dumper_112;
    nodf_module_monitor module_monitor_112;
    nodf_module_intf module_intf_113(clock,reset);
    assign module_intf_113.ap_start = 1'b0;
    assign module_intf_113.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_85_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1226.ap_ready;
    assign module_intf_113.ap_done = 1'b0;
    assign module_intf_113.ap_continue = 1'b0;
    assign module_intf_113.finish = finish;
    csv_file_dump mstatus_csv_dumper_113;
    nodf_module_monitor module_monitor_113;
    nodf_module_intf module_intf_114(clock,reset);
    assign module_intf_114.ap_start = 1'b0;
    assign module_intf_114.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_88_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1234.ap_ready;
    assign module_intf_114.ap_done = 1'b0;
    assign module_intf_114.ap_continue = 1'b0;
    assign module_intf_114.finish = finish;
    csv_file_dump mstatus_csv_dumper_114;
    nodf_module_monitor module_monitor_114;
    nodf_module_intf module_intf_115(clock,reset);
    assign module_intf_115.ap_start = 1'b0;
    assign module_intf_115.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_91_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1243.ap_ready;
    assign module_intf_115.ap_done = 1'b0;
    assign module_intf_115.ap_continue = 1'b0;
    assign module_intf_115.finish = finish;
    csv_file_dump mstatus_csv_dumper_115;
    nodf_module_monitor module_monitor_115;
    nodf_module_intf module_intf_116(clock,reset);
    assign module_intf_116.ap_start = 1'b0;
    assign module_intf_116.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_94_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1252.ap_ready;
    assign module_intf_116.ap_done = 1'b0;
    assign module_intf_116.ap_continue = 1'b0;
    assign module_intf_116.finish = finish;
    csv_file_dump mstatus_csv_dumper_116;
    nodf_module_monitor module_monitor_116;
    nodf_module_intf module_intf_117(clock,reset);
    assign module_intf_117.ap_start = 1'b0;
    assign module_intf_117.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_97_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1261.ap_ready;
    assign module_intf_117.ap_done = 1'b0;
    assign module_intf_117.ap_continue = 1'b0;
    assign module_intf_117.finish = finish;
    csv_file_dump mstatus_csv_dumper_117;
    nodf_module_monitor module_monitor_117;
    nodf_module_intf module_intf_118(clock,reset);
    assign module_intf_118.ap_start = 1'b0;
    assign module_intf_118.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_100_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1270.ap_ready;
    assign module_intf_118.ap_done = 1'b0;
    assign module_intf_118.ap_continue = 1'b0;
    assign module_intf_118.finish = finish;
    csv_file_dump mstatus_csv_dumper_118;
    nodf_module_monitor module_monitor_118;
    nodf_module_intf module_intf_119(clock,reset);
    assign module_intf_119.ap_start = 1'b0;
    assign module_intf_119.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_103_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1278.ap_ready;
    assign module_intf_119.ap_done = 1'b0;
    assign module_intf_119.ap_continue = 1'b0;
    assign module_intf_119.finish = finish;
    csv_file_dump mstatus_csv_dumper_119;
    nodf_module_monitor module_monitor_119;
    nodf_module_intf module_intf_120(clock,reset);
    assign module_intf_120.ap_start = 1'b0;
    assign module_intf_120.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_106_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1287.ap_ready;
    assign module_intf_120.ap_done = 1'b0;
    assign module_intf_120.ap_continue = 1'b0;
    assign module_intf_120.finish = finish;
    csv_file_dump mstatus_csv_dumper_120;
    nodf_module_monitor module_monitor_120;
    nodf_module_intf module_intf_121(clock,reset);
    assign module_intf_121.ap_start = 1'b0;
    assign module_intf_121.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_109_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1296.ap_ready;
    assign module_intf_121.ap_done = 1'b0;
    assign module_intf_121.ap_continue = 1'b0;
    assign module_intf_121.finish = finish;
    csv_file_dump mstatus_csv_dumper_121;
    nodf_module_monitor module_monitor_121;
    nodf_module_intf module_intf_122(clock,reset);
    assign module_intf_122.ap_start = 1'b0;
    assign module_intf_122.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_112_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1305.ap_ready;
    assign module_intf_122.ap_done = 1'b0;
    assign module_intf_122.ap_continue = 1'b0;
    assign module_intf_122.finish = finish;
    csv_file_dump mstatus_csv_dumper_122;
    nodf_module_monitor module_monitor_122;
    nodf_module_intf module_intf_123(clock,reset);
    assign module_intf_123.ap_start = 1'b0;
    assign module_intf_123.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_115_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1314.ap_ready;
    assign module_intf_123.ap_done = 1'b0;
    assign module_intf_123.ap_continue = 1'b0;
    assign module_intf_123.finish = finish;
    csv_file_dump mstatus_csv_dumper_123;
    nodf_module_monitor module_monitor_123;
    nodf_module_intf module_intf_124(clock,reset);
    assign module_intf_124.ap_start = 1'b0;
    assign module_intf_124.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_118_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1322.ap_ready;
    assign module_intf_124.ap_done = 1'b0;
    assign module_intf_124.ap_continue = 1'b0;
    assign module_intf_124.finish = finish;
    csv_file_dump mstatus_csv_dumper_124;
    nodf_module_monitor module_monitor_124;
    nodf_module_intf module_intf_125(clock,reset);
    assign module_intf_125.ap_start = 1'b0;
    assign module_intf_125.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_120_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1331.ap_ready;
    assign module_intf_125.ap_done = 1'b0;
    assign module_intf_125.ap_continue = 1'b0;
    assign module_intf_125.finish = finish;
    csv_file_dump mstatus_csv_dumper_125;
    nodf_module_monitor module_monitor_125;
    nodf_module_intf module_intf_126(clock,reset);
    assign module_intf_126.ap_start = 1'b0;
    assign module_intf_126.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_742.grp_atan2_generic_float_s_fu_169.trunc_ln657_121_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1340.ap_ready;
    assign module_intf_126.ap_done = 1'b0;
    assign module_intf_126.ap_continue = 1'b0;
    assign module_intf_126.finish = finish;
    csv_file_dump mstatus_csv_dumper_126;
    nodf_module_monitor module_monitor_126;
    nodf_module_intf module_intf_127(clock,reset);
    assign module_intf_127.ap_start = 1'b0;
    assign module_intf_127.ap_ready = 1'b0;
    assign module_intf_127.ap_done = 1'b0;
    assign module_intf_127.ap_continue = 1'b0;
    assign module_intf_127.finish = finish;
    csv_file_dump mstatus_csv_dumper_127;
    nodf_module_monitor module_monitor_127;
    nodf_module_intf module_intf_128(clock,reset);
    assign module_intf_128.ap_start = 1'b0;
    assign module_intf_128.ap_ready = 1'b0;
    assign module_intf_128.ap_done = 1'b0;
    assign module_intf_128.ap_continue = 1'b0;
    assign module_intf_128.finish = finish;
    csv_file_dump mstatus_csv_dumper_128;
    nodf_module_monitor module_monitor_128;
    nodf_module_intf module_intf_129(clock,reset);
    assign module_intf_129.ap_start = 1'b0;
    assign module_intf_129.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_8_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_348.ap_ready;
    assign module_intf_129.ap_done = 1'b0;
    assign module_intf_129.ap_continue = 1'b0;
    assign module_intf_129.finish = finish;
    csv_file_dump mstatus_csv_dumper_129;
    nodf_module_monitor module_monitor_129;
    nodf_module_intf module_intf_130(clock,reset);
    assign module_intf_130.ap_start = 1'b0;
    assign module_intf_130.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_1_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_355.ap_ready;
    assign module_intf_130.ap_done = 1'b0;
    assign module_intf_130.ap_continue = 1'b0;
    assign module_intf_130.finish = finish;
    csv_file_dump mstatus_csv_dumper_130;
    nodf_module_monitor module_monitor_130;
    nodf_module_intf module_intf_131(clock,reset);
    assign module_intf_131.ap_start = 1'b0;
    assign module_intf_131.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_4_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_363.ap_ready;
    assign module_intf_131.ap_done = 1'b0;
    assign module_intf_131.ap_continue = 1'b0;
    assign module_intf_131.finish = finish;
    csv_file_dump mstatus_csv_dumper_131;
    nodf_module_monitor module_monitor_131;
    nodf_module_intf module_intf_132(clock,reset);
    assign module_intf_132.ap_start = 1'b0;
    assign module_intf_132.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_7_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_371.ap_ready;
    assign module_intf_132.ap_done = 1'b0;
    assign module_intf_132.ap_continue = 1'b0;
    assign module_intf_132.finish = finish;
    csv_file_dump mstatus_csv_dumper_132;
    nodf_module_monitor module_monitor_132;
    nodf_module_intf module_intf_133(clock,reset);
    assign module_intf_133.ap_start = 1'b0;
    assign module_intf_133.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_12_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_378.ap_ready;
    assign module_intf_133.ap_done = 1'b0;
    assign module_intf_133.ap_continue = 1'b0;
    assign module_intf_133.finish = finish;
    csv_file_dump mstatus_csv_dumper_133;
    nodf_module_monitor module_monitor_133;
    nodf_module_intf module_intf_134(clock,reset);
    assign module_intf_134.ap_start = 1'b0;
    assign module_intf_134.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_15_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_386.ap_ready;
    assign module_intf_134.ap_done = 1'b0;
    assign module_intf_134.ap_continue = 1'b0;
    assign module_intf_134.finish = finish;
    csv_file_dump mstatus_csv_dumper_134;
    nodf_module_monitor module_monitor_134;
    nodf_module_intf module_intf_135(clock,reset);
    assign module_intf_135.ap_start = 1'b0;
    assign module_intf_135.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_18_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_394.ap_ready;
    assign module_intf_135.ap_done = 1'b0;
    assign module_intf_135.ap_continue = 1'b0;
    assign module_intf_135.finish = finish;
    csv_file_dump mstatus_csv_dumper_135;
    nodf_module_monitor module_monitor_135;
    nodf_module_intf module_intf_136(clock,reset);
    assign module_intf_136.ap_start = 1'b0;
    assign module_intf_136.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_21_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_402.ap_ready;
    assign module_intf_136.ap_done = 1'b0;
    assign module_intf_136.ap_continue = 1'b0;
    assign module_intf_136.finish = finish;
    csv_file_dump mstatus_csv_dumper_136;
    nodf_module_monitor module_monitor_136;
    nodf_module_intf module_intf_137(clock,reset);
    assign module_intf_137.ap_start = 1'b0;
    assign module_intf_137.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_24_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_410.ap_ready;
    assign module_intf_137.ap_done = 1'b0;
    assign module_intf_137.ap_continue = 1'b0;
    assign module_intf_137.finish = finish;
    csv_file_dump mstatus_csv_dumper_137;
    nodf_module_monitor module_monitor_137;
    nodf_module_intf module_intf_138(clock,reset);
    assign module_intf_138.ap_start = 1'b0;
    assign module_intf_138.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_27_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_417.ap_ready;
    assign module_intf_138.ap_done = 1'b0;
    assign module_intf_138.ap_continue = 1'b0;
    assign module_intf_138.finish = finish;
    csv_file_dump mstatus_csv_dumper_138;
    nodf_module_monitor module_monitor_138;
    nodf_module_intf module_intf_139(clock,reset);
    assign module_intf_139.ap_start = 1'b0;
    assign module_intf_139.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_30_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_425.ap_ready;
    assign module_intf_139.ap_done = 1'b0;
    assign module_intf_139.ap_continue = 1'b0;
    assign module_intf_139.finish = finish;
    csv_file_dump mstatus_csv_dumper_139;
    nodf_module_monitor module_monitor_139;
    nodf_module_intf module_intf_140(clock,reset);
    assign module_intf_140.ap_start = 1'b0;
    assign module_intf_140.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_33_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_433.ap_ready;
    assign module_intf_140.ap_done = 1'b0;
    assign module_intf_140.ap_continue = 1'b0;
    assign module_intf_140.finish = finish;
    csv_file_dump mstatus_csv_dumper_140;
    nodf_module_monitor module_monitor_140;
    nodf_module_intf module_intf_141(clock,reset);
    assign module_intf_141.ap_start = 1'b0;
    assign module_intf_141.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_36_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_441.ap_ready;
    assign module_intf_141.ap_done = 1'b0;
    assign module_intf_141.ap_continue = 1'b0;
    assign module_intf_141.finish = finish;
    csv_file_dump mstatus_csv_dumper_141;
    nodf_module_monitor module_monitor_141;
    nodf_module_intf module_intf_142(clock,reset);
    assign module_intf_142.ap_start = 1'b0;
    assign module_intf_142.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_39_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_449.ap_ready;
    assign module_intf_142.ap_done = 1'b0;
    assign module_intf_142.ap_continue = 1'b0;
    assign module_intf_142.finish = finish;
    csv_file_dump mstatus_csv_dumper_142;
    nodf_module_monitor module_monitor_142;
    nodf_module_intf module_intf_143(clock,reset);
    assign module_intf_143.ap_start = 1'b0;
    assign module_intf_143.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_42_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_456.ap_ready;
    assign module_intf_143.ap_done = 1'b0;
    assign module_intf_143.ap_continue = 1'b0;
    assign module_intf_143.finish = finish;
    csv_file_dump mstatus_csv_dumper_143;
    nodf_module_monitor module_monitor_143;
    nodf_module_intf module_intf_144(clock,reset);
    assign module_intf_144.ap_start = 1'b0;
    assign module_intf_144.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_45_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_464.ap_ready;
    assign module_intf_144.ap_done = 1'b0;
    assign module_intf_144.ap_continue = 1'b0;
    assign module_intf_144.finish = finish;
    csv_file_dump mstatus_csv_dumper_144;
    nodf_module_monitor module_monitor_144;
    nodf_module_intf module_intf_145(clock,reset);
    assign module_intf_145.ap_start = 1'b0;
    assign module_intf_145.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_48_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_472.ap_ready;
    assign module_intf_145.ap_done = 1'b0;
    assign module_intf_145.ap_continue = 1'b0;
    assign module_intf_145.finish = finish;
    csv_file_dump mstatus_csv_dumper_145;
    nodf_module_monitor module_monitor_145;
    nodf_module_intf module_intf_146(clock,reset);
    assign module_intf_146.ap_start = 1'b0;
    assign module_intf_146.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_51_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_480.ap_ready;
    assign module_intf_146.ap_done = 1'b0;
    assign module_intf_146.ap_continue = 1'b0;
    assign module_intf_146.finish = finish;
    csv_file_dump mstatus_csv_dumper_146;
    nodf_module_monitor module_monitor_146;
    nodf_module_intf module_intf_147(clock,reset);
    assign module_intf_147.ap_start = 1'b0;
    assign module_intf_147.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_54_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_488.ap_ready;
    assign module_intf_147.ap_done = 1'b0;
    assign module_intf_147.ap_continue = 1'b0;
    assign module_intf_147.finish = finish;
    csv_file_dump mstatus_csv_dumper_147;
    nodf_module_monitor module_monitor_147;
    nodf_module_intf module_intf_148(clock,reset);
    assign module_intf_148.ap_start = 1'b0;
    assign module_intf_148.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_57_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_495.ap_ready;
    assign module_intf_148.ap_done = 1'b0;
    assign module_intf_148.ap_continue = 1'b0;
    assign module_intf_148.finish = finish;
    csv_file_dump mstatus_csv_dumper_148;
    nodf_module_monitor module_monitor_148;
    nodf_module_intf module_intf_149(clock,reset);
    assign module_intf_149.ap_start = 1'b0;
    assign module_intf_149.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_60_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_503.ap_ready;
    assign module_intf_149.ap_done = 1'b0;
    assign module_intf_149.ap_continue = 1'b0;
    assign module_intf_149.finish = finish;
    csv_file_dump mstatus_csv_dumper_149;
    nodf_module_monitor module_monitor_149;
    nodf_module_intf module_intf_150(clock,reset);
    assign module_intf_150.ap_start = 1'b0;
    assign module_intf_150.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_63_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_511.ap_ready;
    assign module_intf_150.ap_done = 1'b0;
    assign module_intf_150.ap_continue = 1'b0;
    assign module_intf_150.finish = finish;
    csv_file_dump mstatus_csv_dumper_150;
    nodf_module_monitor module_monitor_150;
    nodf_module_intf module_intf_151(clock,reset);
    assign module_intf_151.ap_start = 1'b0;
    assign module_intf_151.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_66_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_519.ap_ready;
    assign module_intf_151.ap_done = 1'b0;
    assign module_intf_151.ap_continue = 1'b0;
    assign module_intf_151.finish = finish;
    csv_file_dump mstatus_csv_dumper_151;
    nodf_module_monitor module_monitor_151;
    nodf_module_intf module_intf_152(clock,reset);
    assign module_intf_152.ap_start = 1'b0;
    assign module_intf_152.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_69_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_527.ap_ready;
    assign module_intf_152.ap_done = 1'b0;
    assign module_intf_152.ap_continue = 1'b0;
    assign module_intf_152.finish = finish;
    csv_file_dump mstatus_csv_dumper_152;
    nodf_module_monitor module_monitor_152;
    nodf_module_intf module_intf_153(clock,reset);
    assign module_intf_153.ap_start = 1'b0;
    assign module_intf_153.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_72_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_534.ap_ready;
    assign module_intf_153.ap_done = 1'b0;
    assign module_intf_153.ap_continue = 1'b0;
    assign module_intf_153.finish = finish;
    csv_file_dump mstatus_csv_dumper_153;
    nodf_module_monitor module_monitor_153;
    nodf_module_intf module_intf_154(clock,reset);
    assign module_intf_154.ap_start = 1'b0;
    assign module_intf_154.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_75_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_542.ap_ready;
    assign module_intf_154.ap_done = 1'b0;
    assign module_intf_154.ap_continue = 1'b0;
    assign module_intf_154.finish = finish;
    csv_file_dump mstatus_csv_dumper_154;
    nodf_module_monitor module_monitor_154;
    nodf_module_intf module_intf_155(clock,reset);
    assign module_intf_155.ap_start = 1'b0;
    assign module_intf_155.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_78_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_550.ap_ready;
    assign module_intf_155.ap_done = 1'b0;
    assign module_intf_155.ap_continue = 1'b0;
    assign module_intf_155.finish = finish;
    csv_file_dump mstatus_csv_dumper_155;
    nodf_module_monitor module_monitor_155;
    nodf_module_intf module_intf_156(clock,reset);
    assign module_intf_156.ap_start = 1'b0;
    assign module_intf_156.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_81_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_558.ap_ready;
    assign module_intf_156.ap_done = 1'b0;
    assign module_intf_156.ap_continue = 1'b0;
    assign module_intf_156.finish = finish;
    csv_file_dump mstatus_csv_dumper_156;
    nodf_module_monitor module_monitor_156;
    nodf_module_intf module_intf_157(clock,reset);
    assign module_intf_157.ap_start = 1'b0;
    assign module_intf_157.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_84_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_566.ap_ready;
    assign module_intf_157.ap_done = 1'b0;
    assign module_intf_157.ap_continue = 1'b0;
    assign module_intf_157.finish = finish;
    csv_file_dump mstatus_csv_dumper_157;
    nodf_module_monitor module_monitor_157;
    nodf_module_intf module_intf_158(clock,reset);
    assign module_intf_158.ap_start = 1'b0;
    assign module_intf_158.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_87_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_573.ap_ready;
    assign module_intf_158.ap_done = 1'b0;
    assign module_intf_158.ap_continue = 1'b0;
    assign module_intf_158.finish = finish;
    csv_file_dump mstatus_csv_dumper_158;
    nodf_module_monitor module_monitor_158;
    nodf_module_intf module_intf_159(clock,reset);
    assign module_intf_159.ap_start = 1'b0;
    assign module_intf_159.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_90_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_581.ap_ready;
    assign module_intf_159.ap_done = 1'b0;
    assign module_intf_159.ap_continue = 1'b0;
    assign module_intf_159.finish = finish;
    csv_file_dump mstatus_csv_dumper_159;
    nodf_module_monitor module_monitor_159;
    nodf_module_intf module_intf_160(clock,reset);
    assign module_intf_160.ap_start = 1'b0;
    assign module_intf_160.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_93_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_589.ap_ready;
    assign module_intf_160.ap_done = 1'b0;
    assign module_intf_160.ap_continue = 1'b0;
    assign module_intf_160.finish = finish;
    csv_file_dump mstatus_csv_dumper_160;
    nodf_module_monitor module_monitor_160;
    nodf_module_intf module_intf_161(clock,reset);
    assign module_intf_161.ap_start = 1'b0;
    assign module_intf_161.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_96_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_597.ap_ready;
    assign module_intf_161.ap_done = 1'b0;
    assign module_intf_161.ap_continue = 1'b0;
    assign module_intf_161.finish = finish;
    csv_file_dump mstatus_csv_dumper_161;
    nodf_module_monitor module_monitor_161;
    nodf_module_intf module_intf_162(clock,reset);
    assign module_intf_162.ap_start = 1'b0;
    assign module_intf_162.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_99_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_605.ap_ready;
    assign module_intf_162.ap_done = 1'b0;
    assign module_intf_162.ap_continue = 1'b0;
    assign module_intf_162.finish = finish;
    csv_file_dump mstatus_csv_dumper_162;
    nodf_module_monitor module_monitor_162;
    nodf_module_intf module_intf_163(clock,reset);
    assign module_intf_163.ap_start = 1'b0;
    assign module_intf_163.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_102_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_612.ap_ready;
    assign module_intf_163.ap_done = 1'b0;
    assign module_intf_163.ap_continue = 1'b0;
    assign module_intf_163.finish = finish;
    csv_file_dump mstatus_csv_dumper_163;
    nodf_module_monitor module_monitor_163;
    nodf_module_intf module_intf_164(clock,reset);
    assign module_intf_164.ap_start = 1'b0;
    assign module_intf_164.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_105_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_620.ap_ready;
    assign module_intf_164.ap_done = 1'b0;
    assign module_intf_164.ap_continue = 1'b0;
    assign module_intf_164.finish = finish;
    csv_file_dump mstatus_csv_dumper_164;
    nodf_module_monitor module_monitor_164;
    nodf_module_intf module_intf_165(clock,reset);
    assign module_intf_165.ap_start = 1'b0;
    assign module_intf_165.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_108_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_628.ap_ready;
    assign module_intf_165.ap_done = 1'b0;
    assign module_intf_165.ap_continue = 1'b0;
    assign module_intf_165.finish = finish;
    csv_file_dump mstatus_csv_dumper_165;
    nodf_module_monitor module_monitor_165;
    nodf_module_intf module_intf_166(clock,reset);
    assign module_intf_166.ap_start = 1'b0;
    assign module_intf_166.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_111_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_636.ap_ready;
    assign module_intf_166.ap_done = 1'b0;
    assign module_intf_166.ap_continue = 1'b0;
    assign module_intf_166.finish = finish;
    csv_file_dump mstatus_csv_dumper_166;
    nodf_module_monitor module_monitor_166;
    nodf_module_intf module_intf_167(clock,reset);
    assign module_intf_167.ap_start = 1'b0;
    assign module_intf_167.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_114_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_644.ap_ready;
    assign module_intf_167.ap_done = 1'b0;
    assign module_intf_167.ap_continue = 1'b0;
    assign module_intf_167.finish = finish;
    csv_file_dump mstatus_csv_dumper_167;
    nodf_module_monitor module_monitor_167;
    nodf_module_intf module_intf_168(clock,reset);
    assign module_intf_168.ap_start = 1'b0;
    assign module_intf_168.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_117_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_651.ap_ready;
    assign module_intf_168.ap_done = 1'b0;
    assign module_intf_168.ap_continue = 1'b0;
    assign module_intf_168.finish = finish;
    csv_file_dump mstatus_csv_dumper_168;
    nodf_module_monitor module_monitor_168;
    nodf_module_intf module_intf_169(clock,reset);
    assign module_intf_169.ap_start = 1'b0;
    assign module_intf_169.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_119_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_bool_s_fu_659.ap_ready;
    assign module_intf_169.ap_done = 1'b0;
    assign module_intf_169.ap_continue = 1'b0;
    assign module_intf_169.finish = finish;
    csv_file_dump mstatus_csv_dumper_169;
    nodf_module_monitor module_monitor_169;
    nodf_module_intf module_intf_170(clock,reset);
    assign module_intf_170.ap_start = 1'b0;
    assign module_intf_170.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_667.ap_ready;
    assign module_intf_170.ap_done = 1'b0;
    assign module_intf_170.ap_continue = 1'b0;
    assign module_intf_170.finish = finish;
    csv_file_dump mstatus_csv_dumper_170;
    nodf_module_monitor module_monitor_170;
    nodf_module_intf module_intf_171(clock,reset);
    assign module_intf_171.ap_start = 1'b0;
    assign module_intf_171.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_s_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_674.ap_ready;
    assign module_intf_171.ap_done = 1'b0;
    assign module_intf_171.ap_continue = 1'b0;
    assign module_intf_171.finish = finish;
    csv_file_dump mstatus_csv_dumper_171;
    nodf_module_monitor module_monitor_171;
    nodf_module_intf module_intf_172(clock,reset);
    assign module_intf_172.ap_start = 1'b0;
    assign module_intf_172.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_3_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_682.ap_ready;
    assign module_intf_172.ap_done = 1'b0;
    assign module_intf_172.ap_continue = 1'b0;
    assign module_intf_172.finish = finish;
    csv_file_dump mstatus_csv_dumper_172;
    nodf_module_monitor module_monitor_172;
    nodf_module_intf module_intf_173(clock,reset);
    assign module_intf_173.ap_start = 1'b0;
    assign module_intf_173.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_6_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_690.ap_ready;
    assign module_intf_173.ap_done = 1'b0;
    assign module_intf_173.ap_continue = 1'b0;
    assign module_intf_173.finish = finish;
    csv_file_dump mstatus_csv_dumper_173;
    nodf_module_monitor module_monitor_173;
    nodf_module_intf module_intf_174(clock,reset);
    assign module_intf_174.ap_start = 1'b0;
    assign module_intf_174.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_11_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_697.ap_ready;
    assign module_intf_174.ap_done = 1'b0;
    assign module_intf_174.ap_continue = 1'b0;
    assign module_intf_174.finish = finish;
    csv_file_dump mstatus_csv_dumper_174;
    nodf_module_monitor module_monitor_174;
    nodf_module_intf module_intf_175(clock,reset);
    assign module_intf_175.ap_start = 1'b0;
    assign module_intf_175.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_14_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_705.ap_ready;
    assign module_intf_175.ap_done = 1'b0;
    assign module_intf_175.ap_continue = 1'b0;
    assign module_intf_175.finish = finish;
    csv_file_dump mstatus_csv_dumper_175;
    nodf_module_monitor module_monitor_175;
    nodf_module_intf module_intf_176(clock,reset);
    assign module_intf_176.ap_start = 1'b0;
    assign module_intf_176.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_17_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_713.ap_ready;
    assign module_intf_176.ap_done = 1'b0;
    assign module_intf_176.ap_continue = 1'b0;
    assign module_intf_176.finish = finish;
    csv_file_dump mstatus_csv_dumper_176;
    nodf_module_monitor module_monitor_176;
    nodf_module_intf module_intf_177(clock,reset);
    assign module_intf_177.ap_start = 1'b0;
    assign module_intf_177.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_20_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_721.ap_ready;
    assign module_intf_177.ap_done = 1'b0;
    assign module_intf_177.ap_continue = 1'b0;
    assign module_intf_177.finish = finish;
    csv_file_dump mstatus_csv_dumper_177;
    nodf_module_monitor module_monitor_177;
    nodf_module_intf module_intf_178(clock,reset);
    assign module_intf_178.ap_start = 1'b0;
    assign module_intf_178.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_23_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_729.ap_ready;
    assign module_intf_178.ap_done = 1'b0;
    assign module_intf_178.ap_continue = 1'b0;
    assign module_intf_178.finish = finish;
    csv_file_dump mstatus_csv_dumper_178;
    nodf_module_monitor module_monitor_178;
    nodf_module_intf module_intf_179(clock,reset);
    assign module_intf_179.ap_start = 1'b0;
    assign module_intf_179.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_26_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_736.ap_ready;
    assign module_intf_179.ap_done = 1'b0;
    assign module_intf_179.ap_continue = 1'b0;
    assign module_intf_179.finish = finish;
    csv_file_dump mstatus_csv_dumper_179;
    nodf_module_monitor module_monitor_179;
    nodf_module_intf module_intf_180(clock,reset);
    assign module_intf_180.ap_start = 1'b0;
    assign module_intf_180.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_29_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_744.ap_ready;
    assign module_intf_180.ap_done = 1'b0;
    assign module_intf_180.ap_continue = 1'b0;
    assign module_intf_180.finish = finish;
    csv_file_dump mstatus_csv_dumper_180;
    nodf_module_monitor module_monitor_180;
    nodf_module_intf module_intf_181(clock,reset);
    assign module_intf_181.ap_start = 1'b0;
    assign module_intf_181.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_32_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_752.ap_ready;
    assign module_intf_181.ap_done = 1'b0;
    assign module_intf_181.ap_continue = 1'b0;
    assign module_intf_181.finish = finish;
    csv_file_dump mstatus_csv_dumper_181;
    nodf_module_monitor module_monitor_181;
    nodf_module_intf module_intf_182(clock,reset);
    assign module_intf_182.ap_start = 1'b0;
    assign module_intf_182.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_35_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_760.ap_ready;
    assign module_intf_182.ap_done = 1'b0;
    assign module_intf_182.ap_continue = 1'b0;
    assign module_intf_182.finish = finish;
    csv_file_dump mstatus_csv_dumper_182;
    nodf_module_monitor module_monitor_182;
    nodf_module_intf module_intf_183(clock,reset);
    assign module_intf_183.ap_start = 1'b0;
    assign module_intf_183.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_38_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_768.ap_ready;
    assign module_intf_183.ap_done = 1'b0;
    assign module_intf_183.ap_continue = 1'b0;
    assign module_intf_183.finish = finish;
    csv_file_dump mstatus_csv_dumper_183;
    nodf_module_monitor module_monitor_183;
    nodf_module_intf module_intf_184(clock,reset);
    assign module_intf_184.ap_start = 1'b0;
    assign module_intf_184.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_41_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_775.ap_ready;
    assign module_intf_184.ap_done = 1'b0;
    assign module_intf_184.ap_continue = 1'b0;
    assign module_intf_184.finish = finish;
    csv_file_dump mstatus_csv_dumper_184;
    nodf_module_monitor module_monitor_184;
    nodf_module_intf module_intf_185(clock,reset);
    assign module_intf_185.ap_start = 1'b0;
    assign module_intf_185.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_44_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_783.ap_ready;
    assign module_intf_185.ap_done = 1'b0;
    assign module_intf_185.ap_continue = 1'b0;
    assign module_intf_185.finish = finish;
    csv_file_dump mstatus_csv_dumper_185;
    nodf_module_monitor module_monitor_185;
    nodf_module_intf module_intf_186(clock,reset);
    assign module_intf_186.ap_start = 1'b0;
    assign module_intf_186.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_47_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_791.ap_ready;
    assign module_intf_186.ap_done = 1'b0;
    assign module_intf_186.ap_continue = 1'b0;
    assign module_intf_186.finish = finish;
    csv_file_dump mstatus_csv_dumper_186;
    nodf_module_monitor module_monitor_186;
    nodf_module_intf module_intf_187(clock,reset);
    assign module_intf_187.ap_start = 1'b0;
    assign module_intf_187.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_50_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_799.ap_ready;
    assign module_intf_187.ap_done = 1'b0;
    assign module_intf_187.ap_continue = 1'b0;
    assign module_intf_187.finish = finish;
    csv_file_dump mstatus_csv_dumper_187;
    nodf_module_monitor module_monitor_187;
    nodf_module_intf module_intf_188(clock,reset);
    assign module_intf_188.ap_start = 1'b0;
    assign module_intf_188.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_53_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_807.ap_ready;
    assign module_intf_188.ap_done = 1'b0;
    assign module_intf_188.ap_continue = 1'b0;
    assign module_intf_188.finish = finish;
    csv_file_dump mstatus_csv_dumper_188;
    nodf_module_monitor module_monitor_188;
    nodf_module_intf module_intf_189(clock,reset);
    assign module_intf_189.ap_start = 1'b0;
    assign module_intf_189.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_56_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_814.ap_ready;
    assign module_intf_189.ap_done = 1'b0;
    assign module_intf_189.ap_continue = 1'b0;
    assign module_intf_189.finish = finish;
    csv_file_dump mstatus_csv_dumper_189;
    nodf_module_monitor module_monitor_189;
    nodf_module_intf module_intf_190(clock,reset);
    assign module_intf_190.ap_start = 1'b0;
    assign module_intf_190.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_59_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_822.ap_ready;
    assign module_intf_190.ap_done = 1'b0;
    assign module_intf_190.ap_continue = 1'b0;
    assign module_intf_190.finish = finish;
    csv_file_dump mstatus_csv_dumper_190;
    nodf_module_monitor module_monitor_190;
    nodf_module_intf module_intf_191(clock,reset);
    assign module_intf_191.ap_start = 1'b0;
    assign module_intf_191.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_62_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_830.ap_ready;
    assign module_intf_191.ap_done = 1'b0;
    assign module_intf_191.ap_continue = 1'b0;
    assign module_intf_191.finish = finish;
    csv_file_dump mstatus_csv_dumper_191;
    nodf_module_monitor module_monitor_191;
    nodf_module_intf module_intf_192(clock,reset);
    assign module_intf_192.ap_start = 1'b0;
    assign module_intf_192.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_65_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_838.ap_ready;
    assign module_intf_192.ap_done = 1'b0;
    assign module_intf_192.ap_continue = 1'b0;
    assign module_intf_192.finish = finish;
    csv_file_dump mstatus_csv_dumper_192;
    nodf_module_monitor module_monitor_192;
    nodf_module_intf module_intf_193(clock,reset);
    assign module_intf_193.ap_start = 1'b0;
    assign module_intf_193.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_68_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_846.ap_ready;
    assign module_intf_193.ap_done = 1'b0;
    assign module_intf_193.ap_continue = 1'b0;
    assign module_intf_193.finish = finish;
    csv_file_dump mstatus_csv_dumper_193;
    nodf_module_monitor module_monitor_193;
    nodf_module_intf module_intf_194(clock,reset);
    assign module_intf_194.ap_start = 1'b0;
    assign module_intf_194.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_71_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_853.ap_ready;
    assign module_intf_194.ap_done = 1'b0;
    assign module_intf_194.ap_continue = 1'b0;
    assign module_intf_194.finish = finish;
    csv_file_dump mstatus_csv_dumper_194;
    nodf_module_monitor module_monitor_194;
    nodf_module_intf module_intf_195(clock,reset);
    assign module_intf_195.ap_start = 1'b0;
    assign module_intf_195.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_74_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_861.ap_ready;
    assign module_intf_195.ap_done = 1'b0;
    assign module_intf_195.ap_continue = 1'b0;
    assign module_intf_195.finish = finish;
    csv_file_dump mstatus_csv_dumper_195;
    nodf_module_monitor module_monitor_195;
    nodf_module_intf module_intf_196(clock,reset);
    assign module_intf_196.ap_start = 1'b0;
    assign module_intf_196.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_77_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_869.ap_ready;
    assign module_intf_196.ap_done = 1'b0;
    assign module_intf_196.ap_continue = 1'b0;
    assign module_intf_196.finish = finish;
    csv_file_dump mstatus_csv_dumper_196;
    nodf_module_monitor module_monitor_196;
    nodf_module_intf module_intf_197(clock,reset);
    assign module_intf_197.ap_start = 1'b0;
    assign module_intf_197.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_80_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_877.ap_ready;
    assign module_intf_197.ap_done = 1'b0;
    assign module_intf_197.ap_continue = 1'b0;
    assign module_intf_197.finish = finish;
    csv_file_dump mstatus_csv_dumper_197;
    nodf_module_monitor module_monitor_197;
    nodf_module_intf module_intf_198(clock,reset);
    assign module_intf_198.ap_start = 1'b0;
    assign module_intf_198.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_83_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_885.ap_ready;
    assign module_intf_198.ap_done = 1'b0;
    assign module_intf_198.ap_continue = 1'b0;
    assign module_intf_198.finish = finish;
    csv_file_dump mstatus_csv_dumper_198;
    nodf_module_monitor module_monitor_198;
    nodf_module_intf module_intf_199(clock,reset);
    assign module_intf_199.ap_start = 1'b0;
    assign module_intf_199.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_86_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_892.ap_ready;
    assign module_intf_199.ap_done = 1'b0;
    assign module_intf_199.ap_continue = 1'b0;
    assign module_intf_199.finish = finish;
    csv_file_dump mstatus_csv_dumper_199;
    nodf_module_monitor module_monitor_199;
    nodf_module_intf module_intf_200(clock,reset);
    assign module_intf_200.ap_start = 1'b0;
    assign module_intf_200.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_89_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_900.ap_ready;
    assign module_intf_200.ap_done = 1'b0;
    assign module_intf_200.ap_continue = 1'b0;
    assign module_intf_200.finish = finish;
    csv_file_dump mstatus_csv_dumper_200;
    nodf_module_monitor module_monitor_200;
    nodf_module_intf module_intf_201(clock,reset);
    assign module_intf_201.ap_start = 1'b0;
    assign module_intf_201.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_92_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_908.ap_ready;
    assign module_intf_201.ap_done = 1'b0;
    assign module_intf_201.ap_continue = 1'b0;
    assign module_intf_201.finish = finish;
    csv_file_dump mstatus_csv_dumper_201;
    nodf_module_monitor module_monitor_201;
    nodf_module_intf module_intf_202(clock,reset);
    assign module_intf_202.ap_start = 1'b0;
    assign module_intf_202.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_95_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_916.ap_ready;
    assign module_intf_202.ap_done = 1'b0;
    assign module_intf_202.ap_continue = 1'b0;
    assign module_intf_202.finish = finish;
    csv_file_dump mstatus_csv_dumper_202;
    nodf_module_monitor module_monitor_202;
    nodf_module_intf module_intf_203(clock,reset);
    assign module_intf_203.ap_start = 1'b0;
    assign module_intf_203.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_98_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_924.ap_ready;
    assign module_intf_203.ap_done = 1'b0;
    assign module_intf_203.ap_continue = 1'b0;
    assign module_intf_203.finish = finish;
    csv_file_dump mstatus_csv_dumper_203;
    nodf_module_monitor module_monitor_203;
    nodf_module_intf module_intf_204(clock,reset);
    assign module_intf_204.ap_start = 1'b0;
    assign module_intf_204.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_101_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_931.ap_ready;
    assign module_intf_204.ap_done = 1'b0;
    assign module_intf_204.ap_continue = 1'b0;
    assign module_intf_204.finish = finish;
    csv_file_dump mstatus_csv_dumper_204;
    nodf_module_monitor module_monitor_204;
    nodf_module_intf module_intf_205(clock,reset);
    assign module_intf_205.ap_start = 1'b0;
    assign module_intf_205.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_104_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_939.ap_ready;
    assign module_intf_205.ap_done = 1'b0;
    assign module_intf_205.ap_continue = 1'b0;
    assign module_intf_205.finish = finish;
    csv_file_dump mstatus_csv_dumper_205;
    nodf_module_monitor module_monitor_205;
    nodf_module_intf module_intf_206(clock,reset);
    assign module_intf_206.ap_start = 1'b0;
    assign module_intf_206.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_107_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_947.ap_ready;
    assign module_intf_206.ap_done = 1'b0;
    assign module_intf_206.ap_continue = 1'b0;
    assign module_intf_206.finish = finish;
    csv_file_dump mstatus_csv_dumper_206;
    nodf_module_monitor module_monitor_206;
    nodf_module_intf module_intf_207(clock,reset);
    assign module_intf_207.ap_start = 1'b0;
    assign module_intf_207.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_110_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_955.ap_ready;
    assign module_intf_207.ap_done = 1'b0;
    assign module_intf_207.ap_continue = 1'b0;
    assign module_intf_207.finish = finish;
    csv_file_dump mstatus_csv_dumper_207;
    nodf_module_monitor module_monitor_207;
    nodf_module_intf module_intf_208(clock,reset);
    assign module_intf_208.ap_start = 1'b0;
    assign module_intf_208.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_113_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_963.ap_ready;
    assign module_intf_208.ap_done = 1'b0;
    assign module_intf_208.ap_continue = 1'b0;
    assign module_intf_208.finish = finish;
    csv_file_dump mstatus_csv_dumper_208;
    nodf_module_monitor module_monitor_208;
    nodf_module_intf module_intf_209(clock,reset);
    assign module_intf_209.ap_start = 1'b0;
    assign module_intf_209.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_116_addsub_0_0_ap_fixed_43_4_5_3_0_ap_fixed_43_4_5_3_0_ap_uint_1_s_fu_970.ap_ready;
    assign module_intf_209.ap_done = 1'b0;
    assign module_intf_209.ap_continue = 1'b0;
    assign module_intf_209.finish = finish;
    csv_file_dump mstatus_csv_dumper_209;
    nodf_module_monitor module_monitor_209;
    nodf_module_intf module_intf_210(clock,reset);
    assign module_intf_210.ap_start = 1'b0;
    assign module_intf_210.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_9_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_978.ap_ready;
    assign module_intf_210.ap_done = 1'b0;
    assign module_intf_210.ap_continue = 1'b0;
    assign module_intf_210.finish = finish;
    csv_file_dump mstatus_csv_dumper_210;
    nodf_module_monitor module_monitor_210;
    nodf_module_intf module_intf_211(clock,reset);
    assign module_intf_211.ap_start = 1'b0;
    assign module_intf_211.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_2_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_987.ap_ready;
    assign module_intf_211.ap_done = 1'b0;
    assign module_intf_211.ap_continue = 1'b0;
    assign module_intf_211.finish = finish;
    csv_file_dump mstatus_csv_dumper_211;
    nodf_module_monitor module_monitor_211;
    nodf_module_intf module_intf_212(clock,reset);
    assign module_intf_212.ap_start = 1'b0;
    assign module_intf_212.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_5_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_996.ap_ready;
    assign module_intf_212.ap_done = 1'b0;
    assign module_intf_212.ap_continue = 1'b0;
    assign module_intf_212.finish = finish;
    csv_file_dump mstatus_csv_dumper_212;
    nodf_module_monitor module_monitor_212;
    nodf_module_intf module_intf_213(clock,reset);
    assign module_intf_213.ap_start = 1'b0;
    assign module_intf_213.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_10_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1005.ap_ready;
    assign module_intf_213.ap_done = 1'b0;
    assign module_intf_213.ap_continue = 1'b0;
    assign module_intf_213.finish = finish;
    csv_file_dump mstatus_csv_dumper_213;
    nodf_module_monitor module_monitor_213;
    nodf_module_intf module_intf_214(clock,reset);
    assign module_intf_214.ap_start = 1'b0;
    assign module_intf_214.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_13_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1014.ap_ready;
    assign module_intf_214.ap_done = 1'b0;
    assign module_intf_214.ap_continue = 1'b0;
    assign module_intf_214.finish = finish;
    csv_file_dump mstatus_csv_dumper_214;
    nodf_module_monitor module_monitor_214;
    nodf_module_intf module_intf_215(clock,reset);
    assign module_intf_215.ap_start = 1'b0;
    assign module_intf_215.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_16_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1023.ap_ready;
    assign module_intf_215.ap_done = 1'b0;
    assign module_intf_215.ap_continue = 1'b0;
    assign module_intf_215.finish = finish;
    csv_file_dump mstatus_csv_dumper_215;
    nodf_module_monitor module_monitor_215;
    nodf_module_intf module_intf_216(clock,reset);
    assign module_intf_216.ap_start = 1'b0;
    assign module_intf_216.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_19_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1032.ap_ready;
    assign module_intf_216.ap_done = 1'b0;
    assign module_intf_216.ap_continue = 1'b0;
    assign module_intf_216.finish = finish;
    csv_file_dump mstatus_csv_dumper_216;
    nodf_module_monitor module_monitor_216;
    nodf_module_intf module_intf_217(clock,reset);
    assign module_intf_217.ap_start = 1'b0;
    assign module_intf_217.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_22_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1040.ap_ready;
    assign module_intf_217.ap_done = 1'b0;
    assign module_intf_217.ap_continue = 1'b0;
    assign module_intf_217.finish = finish;
    csv_file_dump mstatus_csv_dumper_217;
    nodf_module_monitor module_monitor_217;
    nodf_module_intf module_intf_218(clock,reset);
    assign module_intf_218.ap_start = 1'b0;
    assign module_intf_218.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_25_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1049.ap_ready;
    assign module_intf_218.ap_done = 1'b0;
    assign module_intf_218.ap_continue = 1'b0;
    assign module_intf_218.finish = finish;
    csv_file_dump mstatus_csv_dumper_218;
    nodf_module_monitor module_monitor_218;
    nodf_module_intf module_intf_219(clock,reset);
    assign module_intf_219.ap_start = 1'b0;
    assign module_intf_219.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_28_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1058.ap_ready;
    assign module_intf_219.ap_done = 1'b0;
    assign module_intf_219.ap_continue = 1'b0;
    assign module_intf_219.finish = finish;
    csv_file_dump mstatus_csv_dumper_219;
    nodf_module_monitor module_monitor_219;
    nodf_module_intf module_intf_220(clock,reset);
    assign module_intf_220.ap_start = 1'b0;
    assign module_intf_220.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_31_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1067.ap_ready;
    assign module_intf_220.ap_done = 1'b0;
    assign module_intf_220.ap_continue = 1'b0;
    assign module_intf_220.finish = finish;
    csv_file_dump mstatus_csv_dumper_220;
    nodf_module_monitor module_monitor_220;
    nodf_module_intf module_intf_221(clock,reset);
    assign module_intf_221.ap_start = 1'b0;
    assign module_intf_221.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_34_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1076.ap_ready;
    assign module_intf_221.ap_done = 1'b0;
    assign module_intf_221.ap_continue = 1'b0;
    assign module_intf_221.finish = finish;
    csv_file_dump mstatus_csv_dumper_221;
    nodf_module_monitor module_monitor_221;
    nodf_module_intf module_intf_222(clock,reset);
    assign module_intf_222.ap_start = 1'b0;
    assign module_intf_222.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_37_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1085.ap_ready;
    assign module_intf_222.ap_done = 1'b0;
    assign module_intf_222.ap_continue = 1'b0;
    assign module_intf_222.finish = finish;
    csv_file_dump mstatus_csv_dumper_222;
    nodf_module_monitor module_monitor_222;
    nodf_module_intf module_intf_223(clock,reset);
    assign module_intf_223.ap_start = 1'b0;
    assign module_intf_223.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_40_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1093.ap_ready;
    assign module_intf_223.ap_done = 1'b0;
    assign module_intf_223.ap_continue = 1'b0;
    assign module_intf_223.finish = finish;
    csv_file_dump mstatus_csv_dumper_223;
    nodf_module_monitor module_monitor_223;
    nodf_module_intf module_intf_224(clock,reset);
    assign module_intf_224.ap_start = 1'b0;
    assign module_intf_224.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_43_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1102.ap_ready;
    assign module_intf_224.ap_done = 1'b0;
    assign module_intf_224.ap_continue = 1'b0;
    assign module_intf_224.finish = finish;
    csv_file_dump mstatus_csv_dumper_224;
    nodf_module_monitor module_monitor_224;
    nodf_module_intf module_intf_225(clock,reset);
    assign module_intf_225.ap_start = 1'b0;
    assign module_intf_225.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_46_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1111.ap_ready;
    assign module_intf_225.ap_done = 1'b0;
    assign module_intf_225.ap_continue = 1'b0;
    assign module_intf_225.finish = finish;
    csv_file_dump mstatus_csv_dumper_225;
    nodf_module_monitor module_monitor_225;
    nodf_module_intf module_intf_226(clock,reset);
    assign module_intf_226.ap_start = 1'b0;
    assign module_intf_226.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_49_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1120.ap_ready;
    assign module_intf_226.ap_done = 1'b0;
    assign module_intf_226.ap_continue = 1'b0;
    assign module_intf_226.finish = finish;
    csv_file_dump mstatus_csv_dumper_226;
    nodf_module_monitor module_monitor_226;
    nodf_module_intf module_intf_227(clock,reset);
    assign module_intf_227.ap_start = 1'b0;
    assign module_intf_227.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_52_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1129.ap_ready;
    assign module_intf_227.ap_done = 1'b0;
    assign module_intf_227.ap_continue = 1'b0;
    assign module_intf_227.finish = finish;
    csv_file_dump mstatus_csv_dumper_227;
    nodf_module_monitor module_monitor_227;
    nodf_module_intf module_intf_228(clock,reset);
    assign module_intf_228.ap_start = 1'b0;
    assign module_intf_228.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_55_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1138.ap_ready;
    assign module_intf_228.ap_done = 1'b0;
    assign module_intf_228.ap_continue = 1'b0;
    assign module_intf_228.finish = finish;
    csv_file_dump mstatus_csv_dumper_228;
    nodf_module_monitor module_monitor_228;
    nodf_module_intf module_intf_229(clock,reset);
    assign module_intf_229.ap_start = 1'b0;
    assign module_intf_229.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_58_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1146.ap_ready;
    assign module_intf_229.ap_done = 1'b0;
    assign module_intf_229.ap_continue = 1'b0;
    assign module_intf_229.finish = finish;
    csv_file_dump mstatus_csv_dumper_229;
    nodf_module_monitor module_monitor_229;
    nodf_module_intf module_intf_230(clock,reset);
    assign module_intf_230.ap_start = 1'b0;
    assign module_intf_230.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_61_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1155.ap_ready;
    assign module_intf_230.ap_done = 1'b0;
    assign module_intf_230.ap_continue = 1'b0;
    assign module_intf_230.finish = finish;
    csv_file_dump mstatus_csv_dumper_230;
    nodf_module_monitor module_monitor_230;
    nodf_module_intf module_intf_231(clock,reset);
    assign module_intf_231.ap_start = 1'b0;
    assign module_intf_231.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_64_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1164.ap_ready;
    assign module_intf_231.ap_done = 1'b0;
    assign module_intf_231.ap_continue = 1'b0;
    assign module_intf_231.finish = finish;
    csv_file_dump mstatus_csv_dumper_231;
    nodf_module_monitor module_monitor_231;
    nodf_module_intf module_intf_232(clock,reset);
    assign module_intf_232.ap_start = 1'b0;
    assign module_intf_232.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_67_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1173.ap_ready;
    assign module_intf_232.ap_done = 1'b0;
    assign module_intf_232.ap_continue = 1'b0;
    assign module_intf_232.finish = finish;
    csv_file_dump mstatus_csv_dumper_232;
    nodf_module_monitor module_monitor_232;
    nodf_module_intf module_intf_233(clock,reset);
    assign module_intf_233.ap_start = 1'b0;
    assign module_intf_233.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_70_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1182.ap_ready;
    assign module_intf_233.ap_done = 1'b0;
    assign module_intf_233.ap_continue = 1'b0;
    assign module_intf_233.finish = finish;
    csv_file_dump mstatus_csv_dumper_233;
    nodf_module_monitor module_monitor_233;
    nodf_module_intf module_intf_234(clock,reset);
    assign module_intf_234.ap_start = 1'b0;
    assign module_intf_234.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_73_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1190.ap_ready;
    assign module_intf_234.ap_done = 1'b0;
    assign module_intf_234.ap_continue = 1'b0;
    assign module_intf_234.finish = finish;
    csv_file_dump mstatus_csv_dumper_234;
    nodf_module_monitor module_monitor_234;
    nodf_module_intf module_intf_235(clock,reset);
    assign module_intf_235.ap_start = 1'b0;
    assign module_intf_235.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_76_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1199.ap_ready;
    assign module_intf_235.ap_done = 1'b0;
    assign module_intf_235.ap_continue = 1'b0;
    assign module_intf_235.finish = finish;
    csv_file_dump mstatus_csv_dumper_235;
    nodf_module_monitor module_monitor_235;
    nodf_module_intf module_intf_236(clock,reset);
    assign module_intf_236.ap_start = 1'b0;
    assign module_intf_236.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_79_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1208.ap_ready;
    assign module_intf_236.ap_done = 1'b0;
    assign module_intf_236.ap_continue = 1'b0;
    assign module_intf_236.finish = finish;
    csv_file_dump mstatus_csv_dumper_236;
    nodf_module_monitor module_monitor_236;
    nodf_module_intf module_intf_237(clock,reset);
    assign module_intf_237.ap_start = 1'b0;
    assign module_intf_237.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_82_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1217.ap_ready;
    assign module_intf_237.ap_done = 1'b0;
    assign module_intf_237.ap_continue = 1'b0;
    assign module_intf_237.finish = finish;
    csv_file_dump mstatus_csv_dumper_237;
    nodf_module_monitor module_monitor_237;
    nodf_module_intf module_intf_238(clock,reset);
    assign module_intf_238.ap_start = 1'b0;
    assign module_intf_238.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_85_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1226.ap_ready;
    assign module_intf_238.ap_done = 1'b0;
    assign module_intf_238.ap_continue = 1'b0;
    assign module_intf_238.finish = finish;
    csv_file_dump mstatus_csv_dumper_238;
    nodf_module_monitor module_monitor_238;
    nodf_module_intf module_intf_239(clock,reset);
    assign module_intf_239.ap_start = 1'b0;
    assign module_intf_239.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_88_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1234.ap_ready;
    assign module_intf_239.ap_done = 1'b0;
    assign module_intf_239.ap_continue = 1'b0;
    assign module_intf_239.finish = finish;
    csv_file_dump mstatus_csv_dumper_239;
    nodf_module_monitor module_monitor_239;
    nodf_module_intf module_intf_240(clock,reset);
    assign module_intf_240.ap_start = 1'b0;
    assign module_intf_240.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_91_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1243.ap_ready;
    assign module_intf_240.ap_done = 1'b0;
    assign module_intf_240.ap_continue = 1'b0;
    assign module_intf_240.finish = finish;
    csv_file_dump mstatus_csv_dumper_240;
    nodf_module_monitor module_monitor_240;
    nodf_module_intf module_intf_241(clock,reset);
    assign module_intf_241.ap_start = 1'b0;
    assign module_intf_241.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_94_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1252.ap_ready;
    assign module_intf_241.ap_done = 1'b0;
    assign module_intf_241.ap_continue = 1'b0;
    assign module_intf_241.finish = finish;
    csv_file_dump mstatus_csv_dumper_241;
    nodf_module_monitor module_monitor_241;
    nodf_module_intf module_intf_242(clock,reset);
    assign module_intf_242.ap_start = 1'b0;
    assign module_intf_242.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_97_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1261.ap_ready;
    assign module_intf_242.ap_done = 1'b0;
    assign module_intf_242.ap_continue = 1'b0;
    assign module_intf_242.finish = finish;
    csv_file_dump mstatus_csv_dumper_242;
    nodf_module_monitor module_monitor_242;
    nodf_module_intf module_intf_243(clock,reset);
    assign module_intf_243.ap_start = 1'b0;
    assign module_intf_243.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_100_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1270.ap_ready;
    assign module_intf_243.ap_done = 1'b0;
    assign module_intf_243.ap_continue = 1'b0;
    assign module_intf_243.finish = finish;
    csv_file_dump mstatus_csv_dumper_243;
    nodf_module_monitor module_monitor_243;
    nodf_module_intf module_intf_244(clock,reset);
    assign module_intf_244.ap_start = 1'b0;
    assign module_intf_244.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_103_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1278.ap_ready;
    assign module_intf_244.ap_done = 1'b0;
    assign module_intf_244.ap_continue = 1'b0;
    assign module_intf_244.finish = finish;
    csv_file_dump mstatus_csv_dumper_244;
    nodf_module_monitor module_monitor_244;
    nodf_module_intf module_intf_245(clock,reset);
    assign module_intf_245.ap_start = 1'b0;
    assign module_intf_245.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_106_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1287.ap_ready;
    assign module_intf_245.ap_done = 1'b0;
    assign module_intf_245.ap_continue = 1'b0;
    assign module_intf_245.finish = finish;
    csv_file_dump mstatus_csv_dumper_245;
    nodf_module_monitor module_monitor_245;
    nodf_module_intf module_intf_246(clock,reset);
    assign module_intf_246.ap_start = 1'b0;
    assign module_intf_246.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_109_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1296.ap_ready;
    assign module_intf_246.ap_done = 1'b0;
    assign module_intf_246.ap_continue = 1'b0;
    assign module_intf_246.finish = finish;
    csv_file_dump mstatus_csv_dumper_246;
    nodf_module_monitor module_monitor_246;
    nodf_module_intf module_intf_247(clock,reset);
    assign module_intf_247.ap_start = 1'b0;
    assign module_intf_247.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_112_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1305.ap_ready;
    assign module_intf_247.ap_done = 1'b0;
    assign module_intf_247.ap_continue = 1'b0;
    assign module_intf_247.finish = finish;
    csv_file_dump mstatus_csv_dumper_247;
    nodf_module_monitor module_monitor_247;
    nodf_module_intf module_intf_248(clock,reset);
    assign module_intf_248.ap_start = 1'b0;
    assign module_intf_248.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_115_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1314.ap_ready;
    assign module_intf_248.ap_done = 1'b0;
    assign module_intf_248.ap_continue = 1'b0;
    assign module_intf_248.finish = finish;
    csv_file_dump mstatus_csv_dumper_248;
    nodf_module_monitor module_monitor_248;
    nodf_module_intf module_intf_249(clock,reset);
    assign module_intf_249.ap_start = 1'b0;
    assign module_intf_249.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_118_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1322.ap_ready;
    assign module_intf_249.ap_done = 1'b0;
    assign module_intf_249.ap_continue = 1'b0;
    assign module_intf_249.finish = finish;
    csv_file_dump mstatus_csv_dumper_249;
    nodf_module_monitor module_monitor_249;
    nodf_module_intf module_intf_250(clock,reset);
    assign module_intf_250.ap_start = 1'b0;
    assign module_intf_250.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_120_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1331.ap_ready;
    assign module_intf_250.ap_done = 1'b0;
    assign module_intf_250.ap_continue = 1'b0;
    assign module_intf_250.finish = finish;
    csv_file_dump mstatus_csv_dumper_250;
    nodf_module_monitor module_monitor_250;
    nodf_module_intf module_intf_251(clock,reset);
    assign module_intf_251.ap_start = 1'b0;
    assign module_intf_251.ap_ready = AESL_inst_apskdemod.grp_atan2_cordic_float_s_fu_748.grp_atan2_generic_float_s_fu_169.trunc_ln657_121_addsub_0_0_ap_fixed_40_1_5_3_0_ap_fixed_40_1_0_3_0_ap_uint_1_s_fu_1340.ap_ready;
    assign module_intf_251.ap_done = 1'b0;
    assign module_intf_251.ap_continue = 1'b0;
    assign module_intf_251.finish = finish;
    csv_file_dump mstatus_csv_dumper_251;
    nodf_module_monitor module_monitor_251;
    nodf_module_intf module_intf_252(clock,reset);
    assign module_intf_252.ap_start = AESL_inst_apskdemod.grp_pow_generic_double_s_fu_754.ap_start;
    assign module_intf_252.ap_ready = AESL_inst_apskdemod.grp_pow_generic_double_s_fu_754.ap_ready;
    assign module_intf_252.ap_done = AESL_inst_apskdemod.grp_pow_generic_double_s_fu_754.ap_done;
    assign module_intf_252.ap_continue = 1'b1;
    assign module_intf_252.finish = finish;
    csv_file_dump mstatus_csv_dumper_252;
    nodf_module_monitor module_monitor_252;
    nodf_module_intf module_intf_253(clock,reset);
    assign module_intf_253.ap_start = AESL_inst_apskdemod.grp_pow_generic_double_s_fu_783.ap_start;
    assign module_intf_253.ap_ready = AESL_inst_apskdemod.grp_pow_generic_double_s_fu_783.ap_ready;
    assign module_intf_253.ap_done = AESL_inst_apskdemod.grp_pow_generic_double_s_fu_783.ap_done;
    assign module_intf_253.ap_continue = 1'b1;
    assign module_intf_253.finish = finish;
    csv_file_dump mstatus_csv_dumper_253;
    nodf_module_monitor module_monitor_253;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;



    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);
    mstatus_csv_dumper_5 = new("./module_status5.csv");
    module_monitor_5 = new(module_intf_5,mstatus_csv_dumper_5);
    mstatus_csv_dumper_6 = new("./module_status6.csv");
    module_monitor_6 = new(module_intf_6,mstatus_csv_dumper_6);
    mstatus_csv_dumper_7 = new("./module_status7.csv");
    module_monitor_7 = new(module_intf_7,mstatus_csv_dumper_7);
    mstatus_csv_dumper_8 = new("./module_status8.csv");
    module_monitor_8 = new(module_intf_8,mstatus_csv_dumper_8);
    mstatus_csv_dumper_9 = new("./module_status9.csv");
    module_monitor_9 = new(module_intf_9,mstatus_csv_dumper_9);
    mstatus_csv_dumper_10 = new("./module_status10.csv");
    module_monitor_10 = new(module_intf_10,mstatus_csv_dumper_10);
    mstatus_csv_dumper_11 = new("./module_status11.csv");
    module_monitor_11 = new(module_intf_11,mstatus_csv_dumper_11);
    mstatus_csv_dumper_12 = new("./module_status12.csv");
    module_monitor_12 = new(module_intf_12,mstatus_csv_dumper_12);
    mstatus_csv_dumper_13 = new("./module_status13.csv");
    module_monitor_13 = new(module_intf_13,mstatus_csv_dumper_13);
    mstatus_csv_dumper_14 = new("./module_status14.csv");
    module_monitor_14 = new(module_intf_14,mstatus_csv_dumper_14);
    mstatus_csv_dumper_15 = new("./module_status15.csv");
    module_monitor_15 = new(module_intf_15,mstatus_csv_dumper_15);
    mstatus_csv_dumper_16 = new("./module_status16.csv");
    module_monitor_16 = new(module_intf_16,mstatus_csv_dumper_16);
    mstatus_csv_dumper_17 = new("./module_status17.csv");
    module_monitor_17 = new(module_intf_17,mstatus_csv_dumper_17);
    mstatus_csv_dumper_18 = new("./module_status18.csv");
    module_monitor_18 = new(module_intf_18,mstatus_csv_dumper_18);
    mstatus_csv_dumper_19 = new("./module_status19.csv");
    module_monitor_19 = new(module_intf_19,mstatus_csv_dumper_19);
    mstatus_csv_dumper_20 = new("./module_status20.csv");
    module_monitor_20 = new(module_intf_20,mstatus_csv_dumper_20);
    mstatus_csv_dumper_21 = new("./module_status21.csv");
    module_monitor_21 = new(module_intf_21,mstatus_csv_dumper_21);
    mstatus_csv_dumper_22 = new("./module_status22.csv");
    module_monitor_22 = new(module_intf_22,mstatus_csv_dumper_22);
    mstatus_csv_dumper_23 = new("./module_status23.csv");
    module_monitor_23 = new(module_intf_23,mstatus_csv_dumper_23);
    mstatus_csv_dumper_24 = new("./module_status24.csv");
    module_monitor_24 = new(module_intf_24,mstatus_csv_dumper_24);
    mstatus_csv_dumper_25 = new("./module_status25.csv");
    module_monitor_25 = new(module_intf_25,mstatus_csv_dumper_25);
    mstatus_csv_dumper_26 = new("./module_status26.csv");
    module_monitor_26 = new(module_intf_26,mstatus_csv_dumper_26);
    mstatus_csv_dumper_27 = new("./module_status27.csv");
    module_monitor_27 = new(module_intf_27,mstatus_csv_dumper_27);
    mstatus_csv_dumper_28 = new("./module_status28.csv");
    module_monitor_28 = new(module_intf_28,mstatus_csv_dumper_28);
    mstatus_csv_dumper_29 = new("./module_status29.csv");
    module_monitor_29 = new(module_intf_29,mstatus_csv_dumper_29);
    mstatus_csv_dumper_30 = new("./module_status30.csv");
    module_monitor_30 = new(module_intf_30,mstatus_csv_dumper_30);
    mstatus_csv_dumper_31 = new("./module_status31.csv");
    module_monitor_31 = new(module_intf_31,mstatus_csv_dumper_31);
    mstatus_csv_dumper_32 = new("./module_status32.csv");
    module_monitor_32 = new(module_intf_32,mstatus_csv_dumper_32);
    mstatus_csv_dumper_33 = new("./module_status33.csv");
    module_monitor_33 = new(module_intf_33,mstatus_csv_dumper_33);
    mstatus_csv_dumper_34 = new("./module_status34.csv");
    module_monitor_34 = new(module_intf_34,mstatus_csv_dumper_34);
    mstatus_csv_dumper_35 = new("./module_status35.csv");
    module_monitor_35 = new(module_intf_35,mstatus_csv_dumper_35);
    mstatus_csv_dumper_36 = new("./module_status36.csv");
    module_monitor_36 = new(module_intf_36,mstatus_csv_dumper_36);
    mstatus_csv_dumper_37 = new("./module_status37.csv");
    module_monitor_37 = new(module_intf_37,mstatus_csv_dumper_37);
    mstatus_csv_dumper_38 = new("./module_status38.csv");
    module_monitor_38 = new(module_intf_38,mstatus_csv_dumper_38);
    mstatus_csv_dumper_39 = new("./module_status39.csv");
    module_monitor_39 = new(module_intf_39,mstatus_csv_dumper_39);
    mstatus_csv_dumper_40 = new("./module_status40.csv");
    module_monitor_40 = new(module_intf_40,mstatus_csv_dumper_40);
    mstatus_csv_dumper_41 = new("./module_status41.csv");
    module_monitor_41 = new(module_intf_41,mstatus_csv_dumper_41);
    mstatus_csv_dumper_42 = new("./module_status42.csv");
    module_monitor_42 = new(module_intf_42,mstatus_csv_dumper_42);
    mstatus_csv_dumper_43 = new("./module_status43.csv");
    module_monitor_43 = new(module_intf_43,mstatus_csv_dumper_43);
    mstatus_csv_dumper_44 = new("./module_status44.csv");
    module_monitor_44 = new(module_intf_44,mstatus_csv_dumper_44);
    mstatus_csv_dumper_45 = new("./module_status45.csv");
    module_monitor_45 = new(module_intf_45,mstatus_csv_dumper_45);
    mstatus_csv_dumper_46 = new("./module_status46.csv");
    module_monitor_46 = new(module_intf_46,mstatus_csv_dumper_46);
    mstatus_csv_dumper_47 = new("./module_status47.csv");
    module_monitor_47 = new(module_intf_47,mstatus_csv_dumper_47);
    mstatus_csv_dumper_48 = new("./module_status48.csv");
    module_monitor_48 = new(module_intf_48,mstatus_csv_dumper_48);
    mstatus_csv_dumper_49 = new("./module_status49.csv");
    module_monitor_49 = new(module_intf_49,mstatus_csv_dumper_49);
    mstatus_csv_dumper_50 = new("./module_status50.csv");
    module_monitor_50 = new(module_intf_50,mstatus_csv_dumper_50);
    mstatus_csv_dumper_51 = new("./module_status51.csv");
    module_monitor_51 = new(module_intf_51,mstatus_csv_dumper_51);
    mstatus_csv_dumper_52 = new("./module_status52.csv");
    module_monitor_52 = new(module_intf_52,mstatus_csv_dumper_52);
    mstatus_csv_dumper_53 = new("./module_status53.csv");
    module_monitor_53 = new(module_intf_53,mstatus_csv_dumper_53);
    mstatus_csv_dumper_54 = new("./module_status54.csv");
    module_monitor_54 = new(module_intf_54,mstatus_csv_dumper_54);
    mstatus_csv_dumper_55 = new("./module_status55.csv");
    module_monitor_55 = new(module_intf_55,mstatus_csv_dumper_55);
    mstatus_csv_dumper_56 = new("./module_status56.csv");
    module_monitor_56 = new(module_intf_56,mstatus_csv_dumper_56);
    mstatus_csv_dumper_57 = new("./module_status57.csv");
    module_monitor_57 = new(module_intf_57,mstatus_csv_dumper_57);
    mstatus_csv_dumper_58 = new("./module_status58.csv");
    module_monitor_58 = new(module_intf_58,mstatus_csv_dumper_58);
    mstatus_csv_dumper_59 = new("./module_status59.csv");
    module_monitor_59 = new(module_intf_59,mstatus_csv_dumper_59);
    mstatus_csv_dumper_60 = new("./module_status60.csv");
    module_monitor_60 = new(module_intf_60,mstatus_csv_dumper_60);
    mstatus_csv_dumper_61 = new("./module_status61.csv");
    module_monitor_61 = new(module_intf_61,mstatus_csv_dumper_61);
    mstatus_csv_dumper_62 = new("./module_status62.csv");
    module_monitor_62 = new(module_intf_62,mstatus_csv_dumper_62);
    mstatus_csv_dumper_63 = new("./module_status63.csv");
    module_monitor_63 = new(module_intf_63,mstatus_csv_dumper_63);
    mstatus_csv_dumper_64 = new("./module_status64.csv");
    module_monitor_64 = new(module_intf_64,mstatus_csv_dumper_64);
    mstatus_csv_dumper_65 = new("./module_status65.csv");
    module_monitor_65 = new(module_intf_65,mstatus_csv_dumper_65);
    mstatus_csv_dumper_66 = new("./module_status66.csv");
    module_monitor_66 = new(module_intf_66,mstatus_csv_dumper_66);
    mstatus_csv_dumper_67 = new("./module_status67.csv");
    module_monitor_67 = new(module_intf_67,mstatus_csv_dumper_67);
    mstatus_csv_dumper_68 = new("./module_status68.csv");
    module_monitor_68 = new(module_intf_68,mstatus_csv_dumper_68);
    mstatus_csv_dumper_69 = new("./module_status69.csv");
    module_monitor_69 = new(module_intf_69,mstatus_csv_dumper_69);
    mstatus_csv_dumper_70 = new("./module_status70.csv");
    module_monitor_70 = new(module_intf_70,mstatus_csv_dumper_70);
    mstatus_csv_dumper_71 = new("./module_status71.csv");
    module_monitor_71 = new(module_intf_71,mstatus_csv_dumper_71);
    mstatus_csv_dumper_72 = new("./module_status72.csv");
    module_monitor_72 = new(module_intf_72,mstatus_csv_dumper_72);
    mstatus_csv_dumper_73 = new("./module_status73.csv");
    module_monitor_73 = new(module_intf_73,mstatus_csv_dumper_73);
    mstatus_csv_dumper_74 = new("./module_status74.csv");
    module_monitor_74 = new(module_intf_74,mstatus_csv_dumper_74);
    mstatus_csv_dumper_75 = new("./module_status75.csv");
    module_monitor_75 = new(module_intf_75,mstatus_csv_dumper_75);
    mstatus_csv_dumper_76 = new("./module_status76.csv");
    module_monitor_76 = new(module_intf_76,mstatus_csv_dumper_76);
    mstatus_csv_dumper_77 = new("./module_status77.csv");
    module_monitor_77 = new(module_intf_77,mstatus_csv_dumper_77);
    mstatus_csv_dumper_78 = new("./module_status78.csv");
    module_monitor_78 = new(module_intf_78,mstatus_csv_dumper_78);
    mstatus_csv_dumper_79 = new("./module_status79.csv");
    module_monitor_79 = new(module_intf_79,mstatus_csv_dumper_79);
    mstatus_csv_dumper_80 = new("./module_status80.csv");
    module_monitor_80 = new(module_intf_80,mstatus_csv_dumper_80);
    mstatus_csv_dumper_81 = new("./module_status81.csv");
    module_monitor_81 = new(module_intf_81,mstatus_csv_dumper_81);
    mstatus_csv_dumper_82 = new("./module_status82.csv");
    module_monitor_82 = new(module_intf_82,mstatus_csv_dumper_82);
    mstatus_csv_dumper_83 = new("./module_status83.csv");
    module_monitor_83 = new(module_intf_83,mstatus_csv_dumper_83);
    mstatus_csv_dumper_84 = new("./module_status84.csv");
    module_monitor_84 = new(module_intf_84,mstatus_csv_dumper_84);
    mstatus_csv_dumper_85 = new("./module_status85.csv");
    module_monitor_85 = new(module_intf_85,mstatus_csv_dumper_85);
    mstatus_csv_dumper_86 = new("./module_status86.csv");
    module_monitor_86 = new(module_intf_86,mstatus_csv_dumper_86);
    mstatus_csv_dumper_87 = new("./module_status87.csv");
    module_monitor_87 = new(module_intf_87,mstatus_csv_dumper_87);
    mstatus_csv_dumper_88 = new("./module_status88.csv");
    module_monitor_88 = new(module_intf_88,mstatus_csv_dumper_88);
    mstatus_csv_dumper_89 = new("./module_status89.csv");
    module_monitor_89 = new(module_intf_89,mstatus_csv_dumper_89);
    mstatus_csv_dumper_90 = new("./module_status90.csv");
    module_monitor_90 = new(module_intf_90,mstatus_csv_dumper_90);
    mstatus_csv_dumper_91 = new("./module_status91.csv");
    module_monitor_91 = new(module_intf_91,mstatus_csv_dumper_91);
    mstatus_csv_dumper_92 = new("./module_status92.csv");
    module_monitor_92 = new(module_intf_92,mstatus_csv_dumper_92);
    mstatus_csv_dumper_93 = new("./module_status93.csv");
    module_monitor_93 = new(module_intf_93,mstatus_csv_dumper_93);
    mstatus_csv_dumper_94 = new("./module_status94.csv");
    module_monitor_94 = new(module_intf_94,mstatus_csv_dumper_94);
    mstatus_csv_dumper_95 = new("./module_status95.csv");
    module_monitor_95 = new(module_intf_95,mstatus_csv_dumper_95);
    mstatus_csv_dumper_96 = new("./module_status96.csv");
    module_monitor_96 = new(module_intf_96,mstatus_csv_dumper_96);
    mstatus_csv_dumper_97 = new("./module_status97.csv");
    module_monitor_97 = new(module_intf_97,mstatus_csv_dumper_97);
    mstatus_csv_dumper_98 = new("./module_status98.csv");
    module_monitor_98 = new(module_intf_98,mstatus_csv_dumper_98);
    mstatus_csv_dumper_99 = new("./module_status99.csv");
    module_monitor_99 = new(module_intf_99,mstatus_csv_dumper_99);
    mstatus_csv_dumper_100 = new("./module_status100.csv");
    module_monitor_100 = new(module_intf_100,mstatus_csv_dumper_100);
    mstatus_csv_dumper_101 = new("./module_status101.csv");
    module_monitor_101 = new(module_intf_101,mstatus_csv_dumper_101);
    mstatus_csv_dumper_102 = new("./module_status102.csv");
    module_monitor_102 = new(module_intf_102,mstatus_csv_dumper_102);
    mstatus_csv_dumper_103 = new("./module_status103.csv");
    module_monitor_103 = new(module_intf_103,mstatus_csv_dumper_103);
    mstatus_csv_dumper_104 = new("./module_status104.csv");
    module_monitor_104 = new(module_intf_104,mstatus_csv_dumper_104);
    mstatus_csv_dumper_105 = new("./module_status105.csv");
    module_monitor_105 = new(module_intf_105,mstatus_csv_dumper_105);
    mstatus_csv_dumper_106 = new("./module_status106.csv");
    module_monitor_106 = new(module_intf_106,mstatus_csv_dumper_106);
    mstatus_csv_dumper_107 = new("./module_status107.csv");
    module_monitor_107 = new(module_intf_107,mstatus_csv_dumper_107);
    mstatus_csv_dumper_108 = new("./module_status108.csv");
    module_monitor_108 = new(module_intf_108,mstatus_csv_dumper_108);
    mstatus_csv_dumper_109 = new("./module_status109.csv");
    module_monitor_109 = new(module_intf_109,mstatus_csv_dumper_109);
    mstatus_csv_dumper_110 = new("./module_status110.csv");
    module_monitor_110 = new(module_intf_110,mstatus_csv_dumper_110);
    mstatus_csv_dumper_111 = new("./module_status111.csv");
    module_monitor_111 = new(module_intf_111,mstatus_csv_dumper_111);
    mstatus_csv_dumper_112 = new("./module_status112.csv");
    module_monitor_112 = new(module_intf_112,mstatus_csv_dumper_112);
    mstatus_csv_dumper_113 = new("./module_status113.csv");
    module_monitor_113 = new(module_intf_113,mstatus_csv_dumper_113);
    mstatus_csv_dumper_114 = new("./module_status114.csv");
    module_monitor_114 = new(module_intf_114,mstatus_csv_dumper_114);
    mstatus_csv_dumper_115 = new("./module_status115.csv");
    module_monitor_115 = new(module_intf_115,mstatus_csv_dumper_115);
    mstatus_csv_dumper_116 = new("./module_status116.csv");
    module_monitor_116 = new(module_intf_116,mstatus_csv_dumper_116);
    mstatus_csv_dumper_117 = new("./module_status117.csv");
    module_monitor_117 = new(module_intf_117,mstatus_csv_dumper_117);
    mstatus_csv_dumper_118 = new("./module_status118.csv");
    module_monitor_118 = new(module_intf_118,mstatus_csv_dumper_118);
    mstatus_csv_dumper_119 = new("./module_status119.csv");
    module_monitor_119 = new(module_intf_119,mstatus_csv_dumper_119);
    mstatus_csv_dumper_120 = new("./module_status120.csv");
    module_monitor_120 = new(module_intf_120,mstatus_csv_dumper_120);
    mstatus_csv_dumper_121 = new("./module_status121.csv");
    module_monitor_121 = new(module_intf_121,mstatus_csv_dumper_121);
    mstatus_csv_dumper_122 = new("./module_status122.csv");
    module_monitor_122 = new(module_intf_122,mstatus_csv_dumper_122);
    mstatus_csv_dumper_123 = new("./module_status123.csv");
    module_monitor_123 = new(module_intf_123,mstatus_csv_dumper_123);
    mstatus_csv_dumper_124 = new("./module_status124.csv");
    module_monitor_124 = new(module_intf_124,mstatus_csv_dumper_124);
    mstatus_csv_dumper_125 = new("./module_status125.csv");
    module_monitor_125 = new(module_intf_125,mstatus_csv_dumper_125);
    mstatus_csv_dumper_126 = new("./module_status126.csv");
    module_monitor_126 = new(module_intf_126,mstatus_csv_dumper_126);
    mstatus_csv_dumper_127 = new("./module_status127.csv");
    module_monitor_127 = new(module_intf_127,mstatus_csv_dumper_127);
    mstatus_csv_dumper_128 = new("./module_status128.csv");
    module_monitor_128 = new(module_intf_128,mstatus_csv_dumper_128);
    mstatus_csv_dumper_129 = new("./module_status129.csv");
    module_monitor_129 = new(module_intf_129,mstatus_csv_dumper_129);
    mstatus_csv_dumper_130 = new("./module_status130.csv");
    module_monitor_130 = new(module_intf_130,mstatus_csv_dumper_130);
    mstatus_csv_dumper_131 = new("./module_status131.csv");
    module_monitor_131 = new(module_intf_131,mstatus_csv_dumper_131);
    mstatus_csv_dumper_132 = new("./module_status132.csv");
    module_monitor_132 = new(module_intf_132,mstatus_csv_dumper_132);
    mstatus_csv_dumper_133 = new("./module_status133.csv");
    module_monitor_133 = new(module_intf_133,mstatus_csv_dumper_133);
    mstatus_csv_dumper_134 = new("./module_status134.csv");
    module_monitor_134 = new(module_intf_134,mstatus_csv_dumper_134);
    mstatus_csv_dumper_135 = new("./module_status135.csv");
    module_monitor_135 = new(module_intf_135,mstatus_csv_dumper_135);
    mstatus_csv_dumper_136 = new("./module_status136.csv");
    module_monitor_136 = new(module_intf_136,mstatus_csv_dumper_136);
    mstatus_csv_dumper_137 = new("./module_status137.csv");
    module_monitor_137 = new(module_intf_137,mstatus_csv_dumper_137);
    mstatus_csv_dumper_138 = new("./module_status138.csv");
    module_monitor_138 = new(module_intf_138,mstatus_csv_dumper_138);
    mstatus_csv_dumper_139 = new("./module_status139.csv");
    module_monitor_139 = new(module_intf_139,mstatus_csv_dumper_139);
    mstatus_csv_dumper_140 = new("./module_status140.csv");
    module_monitor_140 = new(module_intf_140,mstatus_csv_dumper_140);
    mstatus_csv_dumper_141 = new("./module_status141.csv");
    module_monitor_141 = new(module_intf_141,mstatus_csv_dumper_141);
    mstatus_csv_dumper_142 = new("./module_status142.csv");
    module_monitor_142 = new(module_intf_142,mstatus_csv_dumper_142);
    mstatus_csv_dumper_143 = new("./module_status143.csv");
    module_monitor_143 = new(module_intf_143,mstatus_csv_dumper_143);
    mstatus_csv_dumper_144 = new("./module_status144.csv");
    module_monitor_144 = new(module_intf_144,mstatus_csv_dumper_144);
    mstatus_csv_dumper_145 = new("./module_status145.csv");
    module_monitor_145 = new(module_intf_145,mstatus_csv_dumper_145);
    mstatus_csv_dumper_146 = new("./module_status146.csv");
    module_monitor_146 = new(module_intf_146,mstatus_csv_dumper_146);
    mstatus_csv_dumper_147 = new("./module_status147.csv");
    module_monitor_147 = new(module_intf_147,mstatus_csv_dumper_147);
    mstatus_csv_dumper_148 = new("./module_status148.csv");
    module_monitor_148 = new(module_intf_148,mstatus_csv_dumper_148);
    mstatus_csv_dumper_149 = new("./module_status149.csv");
    module_monitor_149 = new(module_intf_149,mstatus_csv_dumper_149);
    mstatus_csv_dumper_150 = new("./module_status150.csv");
    module_monitor_150 = new(module_intf_150,mstatus_csv_dumper_150);
    mstatus_csv_dumper_151 = new("./module_status151.csv");
    module_monitor_151 = new(module_intf_151,mstatus_csv_dumper_151);
    mstatus_csv_dumper_152 = new("./module_status152.csv");
    module_monitor_152 = new(module_intf_152,mstatus_csv_dumper_152);
    mstatus_csv_dumper_153 = new("./module_status153.csv");
    module_monitor_153 = new(module_intf_153,mstatus_csv_dumper_153);
    mstatus_csv_dumper_154 = new("./module_status154.csv");
    module_monitor_154 = new(module_intf_154,mstatus_csv_dumper_154);
    mstatus_csv_dumper_155 = new("./module_status155.csv");
    module_monitor_155 = new(module_intf_155,mstatus_csv_dumper_155);
    mstatus_csv_dumper_156 = new("./module_status156.csv");
    module_monitor_156 = new(module_intf_156,mstatus_csv_dumper_156);
    mstatus_csv_dumper_157 = new("./module_status157.csv");
    module_monitor_157 = new(module_intf_157,mstatus_csv_dumper_157);
    mstatus_csv_dumper_158 = new("./module_status158.csv");
    module_monitor_158 = new(module_intf_158,mstatus_csv_dumper_158);
    mstatus_csv_dumper_159 = new("./module_status159.csv");
    module_monitor_159 = new(module_intf_159,mstatus_csv_dumper_159);
    mstatus_csv_dumper_160 = new("./module_status160.csv");
    module_monitor_160 = new(module_intf_160,mstatus_csv_dumper_160);
    mstatus_csv_dumper_161 = new("./module_status161.csv");
    module_monitor_161 = new(module_intf_161,mstatus_csv_dumper_161);
    mstatus_csv_dumper_162 = new("./module_status162.csv");
    module_monitor_162 = new(module_intf_162,mstatus_csv_dumper_162);
    mstatus_csv_dumper_163 = new("./module_status163.csv");
    module_monitor_163 = new(module_intf_163,mstatus_csv_dumper_163);
    mstatus_csv_dumper_164 = new("./module_status164.csv");
    module_monitor_164 = new(module_intf_164,mstatus_csv_dumper_164);
    mstatus_csv_dumper_165 = new("./module_status165.csv");
    module_monitor_165 = new(module_intf_165,mstatus_csv_dumper_165);
    mstatus_csv_dumper_166 = new("./module_status166.csv");
    module_monitor_166 = new(module_intf_166,mstatus_csv_dumper_166);
    mstatus_csv_dumper_167 = new("./module_status167.csv");
    module_monitor_167 = new(module_intf_167,mstatus_csv_dumper_167);
    mstatus_csv_dumper_168 = new("./module_status168.csv");
    module_monitor_168 = new(module_intf_168,mstatus_csv_dumper_168);
    mstatus_csv_dumper_169 = new("./module_status169.csv");
    module_monitor_169 = new(module_intf_169,mstatus_csv_dumper_169);
    mstatus_csv_dumper_170 = new("./module_status170.csv");
    module_monitor_170 = new(module_intf_170,mstatus_csv_dumper_170);
    mstatus_csv_dumper_171 = new("./module_status171.csv");
    module_monitor_171 = new(module_intf_171,mstatus_csv_dumper_171);
    mstatus_csv_dumper_172 = new("./module_status172.csv");
    module_monitor_172 = new(module_intf_172,mstatus_csv_dumper_172);
    mstatus_csv_dumper_173 = new("./module_status173.csv");
    module_monitor_173 = new(module_intf_173,mstatus_csv_dumper_173);
    mstatus_csv_dumper_174 = new("./module_status174.csv");
    module_monitor_174 = new(module_intf_174,mstatus_csv_dumper_174);
    mstatus_csv_dumper_175 = new("./module_status175.csv");
    module_monitor_175 = new(module_intf_175,mstatus_csv_dumper_175);
    mstatus_csv_dumper_176 = new("./module_status176.csv");
    module_monitor_176 = new(module_intf_176,mstatus_csv_dumper_176);
    mstatus_csv_dumper_177 = new("./module_status177.csv");
    module_monitor_177 = new(module_intf_177,mstatus_csv_dumper_177);
    mstatus_csv_dumper_178 = new("./module_status178.csv");
    module_monitor_178 = new(module_intf_178,mstatus_csv_dumper_178);
    mstatus_csv_dumper_179 = new("./module_status179.csv");
    module_monitor_179 = new(module_intf_179,mstatus_csv_dumper_179);
    mstatus_csv_dumper_180 = new("./module_status180.csv");
    module_monitor_180 = new(module_intf_180,mstatus_csv_dumper_180);
    mstatus_csv_dumper_181 = new("./module_status181.csv");
    module_monitor_181 = new(module_intf_181,mstatus_csv_dumper_181);
    mstatus_csv_dumper_182 = new("./module_status182.csv");
    module_monitor_182 = new(module_intf_182,mstatus_csv_dumper_182);
    mstatus_csv_dumper_183 = new("./module_status183.csv");
    module_monitor_183 = new(module_intf_183,mstatus_csv_dumper_183);
    mstatus_csv_dumper_184 = new("./module_status184.csv");
    module_monitor_184 = new(module_intf_184,mstatus_csv_dumper_184);
    mstatus_csv_dumper_185 = new("./module_status185.csv");
    module_monitor_185 = new(module_intf_185,mstatus_csv_dumper_185);
    mstatus_csv_dumper_186 = new("./module_status186.csv");
    module_monitor_186 = new(module_intf_186,mstatus_csv_dumper_186);
    mstatus_csv_dumper_187 = new("./module_status187.csv");
    module_monitor_187 = new(module_intf_187,mstatus_csv_dumper_187);
    mstatus_csv_dumper_188 = new("./module_status188.csv");
    module_monitor_188 = new(module_intf_188,mstatus_csv_dumper_188);
    mstatus_csv_dumper_189 = new("./module_status189.csv");
    module_monitor_189 = new(module_intf_189,mstatus_csv_dumper_189);
    mstatus_csv_dumper_190 = new("./module_status190.csv");
    module_monitor_190 = new(module_intf_190,mstatus_csv_dumper_190);
    mstatus_csv_dumper_191 = new("./module_status191.csv");
    module_monitor_191 = new(module_intf_191,mstatus_csv_dumper_191);
    mstatus_csv_dumper_192 = new("./module_status192.csv");
    module_monitor_192 = new(module_intf_192,mstatus_csv_dumper_192);
    mstatus_csv_dumper_193 = new("./module_status193.csv");
    module_monitor_193 = new(module_intf_193,mstatus_csv_dumper_193);
    mstatus_csv_dumper_194 = new("./module_status194.csv");
    module_monitor_194 = new(module_intf_194,mstatus_csv_dumper_194);
    mstatus_csv_dumper_195 = new("./module_status195.csv");
    module_monitor_195 = new(module_intf_195,mstatus_csv_dumper_195);
    mstatus_csv_dumper_196 = new("./module_status196.csv");
    module_monitor_196 = new(module_intf_196,mstatus_csv_dumper_196);
    mstatus_csv_dumper_197 = new("./module_status197.csv");
    module_monitor_197 = new(module_intf_197,mstatus_csv_dumper_197);
    mstatus_csv_dumper_198 = new("./module_status198.csv");
    module_monitor_198 = new(module_intf_198,mstatus_csv_dumper_198);
    mstatus_csv_dumper_199 = new("./module_status199.csv");
    module_monitor_199 = new(module_intf_199,mstatus_csv_dumper_199);
    mstatus_csv_dumper_200 = new("./module_status200.csv");
    module_monitor_200 = new(module_intf_200,mstatus_csv_dumper_200);
    mstatus_csv_dumper_201 = new("./module_status201.csv");
    module_monitor_201 = new(module_intf_201,mstatus_csv_dumper_201);
    mstatus_csv_dumper_202 = new("./module_status202.csv");
    module_monitor_202 = new(module_intf_202,mstatus_csv_dumper_202);
    mstatus_csv_dumper_203 = new("./module_status203.csv");
    module_monitor_203 = new(module_intf_203,mstatus_csv_dumper_203);
    mstatus_csv_dumper_204 = new("./module_status204.csv");
    module_monitor_204 = new(module_intf_204,mstatus_csv_dumper_204);
    mstatus_csv_dumper_205 = new("./module_status205.csv");
    module_monitor_205 = new(module_intf_205,mstatus_csv_dumper_205);
    mstatus_csv_dumper_206 = new("./module_status206.csv");
    module_monitor_206 = new(module_intf_206,mstatus_csv_dumper_206);
    mstatus_csv_dumper_207 = new("./module_status207.csv");
    module_monitor_207 = new(module_intf_207,mstatus_csv_dumper_207);
    mstatus_csv_dumper_208 = new("./module_status208.csv");
    module_monitor_208 = new(module_intf_208,mstatus_csv_dumper_208);
    mstatus_csv_dumper_209 = new("./module_status209.csv");
    module_monitor_209 = new(module_intf_209,mstatus_csv_dumper_209);
    mstatus_csv_dumper_210 = new("./module_status210.csv");
    module_monitor_210 = new(module_intf_210,mstatus_csv_dumper_210);
    mstatus_csv_dumper_211 = new("./module_status211.csv");
    module_monitor_211 = new(module_intf_211,mstatus_csv_dumper_211);
    mstatus_csv_dumper_212 = new("./module_status212.csv");
    module_monitor_212 = new(module_intf_212,mstatus_csv_dumper_212);
    mstatus_csv_dumper_213 = new("./module_status213.csv");
    module_monitor_213 = new(module_intf_213,mstatus_csv_dumper_213);
    mstatus_csv_dumper_214 = new("./module_status214.csv");
    module_monitor_214 = new(module_intf_214,mstatus_csv_dumper_214);
    mstatus_csv_dumper_215 = new("./module_status215.csv");
    module_monitor_215 = new(module_intf_215,mstatus_csv_dumper_215);
    mstatus_csv_dumper_216 = new("./module_status216.csv");
    module_monitor_216 = new(module_intf_216,mstatus_csv_dumper_216);
    mstatus_csv_dumper_217 = new("./module_status217.csv");
    module_monitor_217 = new(module_intf_217,mstatus_csv_dumper_217);
    mstatus_csv_dumper_218 = new("./module_status218.csv");
    module_monitor_218 = new(module_intf_218,mstatus_csv_dumper_218);
    mstatus_csv_dumper_219 = new("./module_status219.csv");
    module_monitor_219 = new(module_intf_219,mstatus_csv_dumper_219);
    mstatus_csv_dumper_220 = new("./module_status220.csv");
    module_monitor_220 = new(module_intf_220,mstatus_csv_dumper_220);
    mstatus_csv_dumper_221 = new("./module_status221.csv");
    module_monitor_221 = new(module_intf_221,mstatus_csv_dumper_221);
    mstatus_csv_dumper_222 = new("./module_status222.csv");
    module_monitor_222 = new(module_intf_222,mstatus_csv_dumper_222);
    mstatus_csv_dumper_223 = new("./module_status223.csv");
    module_monitor_223 = new(module_intf_223,mstatus_csv_dumper_223);
    mstatus_csv_dumper_224 = new("./module_status224.csv");
    module_monitor_224 = new(module_intf_224,mstatus_csv_dumper_224);
    mstatus_csv_dumper_225 = new("./module_status225.csv");
    module_monitor_225 = new(module_intf_225,mstatus_csv_dumper_225);
    mstatus_csv_dumper_226 = new("./module_status226.csv");
    module_monitor_226 = new(module_intf_226,mstatus_csv_dumper_226);
    mstatus_csv_dumper_227 = new("./module_status227.csv");
    module_monitor_227 = new(module_intf_227,mstatus_csv_dumper_227);
    mstatus_csv_dumper_228 = new("./module_status228.csv");
    module_monitor_228 = new(module_intf_228,mstatus_csv_dumper_228);
    mstatus_csv_dumper_229 = new("./module_status229.csv");
    module_monitor_229 = new(module_intf_229,mstatus_csv_dumper_229);
    mstatus_csv_dumper_230 = new("./module_status230.csv");
    module_monitor_230 = new(module_intf_230,mstatus_csv_dumper_230);
    mstatus_csv_dumper_231 = new("./module_status231.csv");
    module_monitor_231 = new(module_intf_231,mstatus_csv_dumper_231);
    mstatus_csv_dumper_232 = new("./module_status232.csv");
    module_monitor_232 = new(module_intf_232,mstatus_csv_dumper_232);
    mstatus_csv_dumper_233 = new("./module_status233.csv");
    module_monitor_233 = new(module_intf_233,mstatus_csv_dumper_233);
    mstatus_csv_dumper_234 = new("./module_status234.csv");
    module_monitor_234 = new(module_intf_234,mstatus_csv_dumper_234);
    mstatus_csv_dumper_235 = new("./module_status235.csv");
    module_monitor_235 = new(module_intf_235,mstatus_csv_dumper_235);
    mstatus_csv_dumper_236 = new("./module_status236.csv");
    module_monitor_236 = new(module_intf_236,mstatus_csv_dumper_236);
    mstatus_csv_dumper_237 = new("./module_status237.csv");
    module_monitor_237 = new(module_intf_237,mstatus_csv_dumper_237);
    mstatus_csv_dumper_238 = new("./module_status238.csv");
    module_monitor_238 = new(module_intf_238,mstatus_csv_dumper_238);
    mstatus_csv_dumper_239 = new("./module_status239.csv");
    module_monitor_239 = new(module_intf_239,mstatus_csv_dumper_239);
    mstatus_csv_dumper_240 = new("./module_status240.csv");
    module_monitor_240 = new(module_intf_240,mstatus_csv_dumper_240);
    mstatus_csv_dumper_241 = new("./module_status241.csv");
    module_monitor_241 = new(module_intf_241,mstatus_csv_dumper_241);
    mstatus_csv_dumper_242 = new("./module_status242.csv");
    module_monitor_242 = new(module_intf_242,mstatus_csv_dumper_242);
    mstatus_csv_dumper_243 = new("./module_status243.csv");
    module_monitor_243 = new(module_intf_243,mstatus_csv_dumper_243);
    mstatus_csv_dumper_244 = new("./module_status244.csv");
    module_monitor_244 = new(module_intf_244,mstatus_csv_dumper_244);
    mstatus_csv_dumper_245 = new("./module_status245.csv");
    module_monitor_245 = new(module_intf_245,mstatus_csv_dumper_245);
    mstatus_csv_dumper_246 = new("./module_status246.csv");
    module_monitor_246 = new(module_intf_246,mstatus_csv_dumper_246);
    mstatus_csv_dumper_247 = new("./module_status247.csv");
    module_monitor_247 = new(module_intf_247,mstatus_csv_dumper_247);
    mstatus_csv_dumper_248 = new("./module_status248.csv");
    module_monitor_248 = new(module_intf_248,mstatus_csv_dumper_248);
    mstatus_csv_dumper_249 = new("./module_status249.csv");
    module_monitor_249 = new(module_intf_249,mstatus_csv_dumper_249);
    mstatus_csv_dumper_250 = new("./module_status250.csv");
    module_monitor_250 = new(module_intf_250,mstatus_csv_dumper_250);
    mstatus_csv_dumper_251 = new("./module_status251.csv");
    module_monitor_251 = new(module_intf_251,mstatus_csv_dumper_251);
    mstatus_csv_dumper_252 = new("./module_status252.csv");
    module_monitor_252 = new(module_intf_252,mstatus_csv_dumper_252);
    mstatus_csv_dumper_253 = new("./module_status253.csv");
    module_monitor_253 = new(module_intf_253,mstatus_csv_dumper_253);

    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_6);
    sample_manager_inst.add_one_monitor(module_monitor_7);
    sample_manager_inst.add_one_monitor(module_monitor_8);
    sample_manager_inst.add_one_monitor(module_monitor_9);
    sample_manager_inst.add_one_monitor(module_monitor_10);
    sample_manager_inst.add_one_monitor(module_monitor_11);
    sample_manager_inst.add_one_monitor(module_monitor_12);
    sample_manager_inst.add_one_monitor(module_monitor_13);
    sample_manager_inst.add_one_monitor(module_monitor_14);
    sample_manager_inst.add_one_monitor(module_monitor_15);
    sample_manager_inst.add_one_monitor(module_monitor_16);
    sample_manager_inst.add_one_monitor(module_monitor_17);
    sample_manager_inst.add_one_monitor(module_monitor_18);
    sample_manager_inst.add_one_monitor(module_monitor_19);
    sample_manager_inst.add_one_monitor(module_monitor_20);
    sample_manager_inst.add_one_monitor(module_monitor_21);
    sample_manager_inst.add_one_monitor(module_monitor_22);
    sample_manager_inst.add_one_monitor(module_monitor_23);
    sample_manager_inst.add_one_monitor(module_monitor_24);
    sample_manager_inst.add_one_monitor(module_monitor_25);
    sample_manager_inst.add_one_monitor(module_monitor_26);
    sample_manager_inst.add_one_monitor(module_monitor_27);
    sample_manager_inst.add_one_monitor(module_monitor_28);
    sample_manager_inst.add_one_monitor(module_monitor_29);
    sample_manager_inst.add_one_monitor(module_monitor_30);
    sample_manager_inst.add_one_monitor(module_monitor_31);
    sample_manager_inst.add_one_monitor(module_monitor_32);
    sample_manager_inst.add_one_monitor(module_monitor_33);
    sample_manager_inst.add_one_monitor(module_monitor_34);
    sample_manager_inst.add_one_monitor(module_monitor_35);
    sample_manager_inst.add_one_monitor(module_monitor_36);
    sample_manager_inst.add_one_monitor(module_monitor_37);
    sample_manager_inst.add_one_monitor(module_monitor_38);
    sample_manager_inst.add_one_monitor(module_monitor_39);
    sample_manager_inst.add_one_monitor(module_monitor_40);
    sample_manager_inst.add_one_monitor(module_monitor_41);
    sample_manager_inst.add_one_monitor(module_monitor_42);
    sample_manager_inst.add_one_monitor(module_monitor_43);
    sample_manager_inst.add_one_monitor(module_monitor_44);
    sample_manager_inst.add_one_monitor(module_monitor_45);
    sample_manager_inst.add_one_monitor(module_monitor_46);
    sample_manager_inst.add_one_monitor(module_monitor_47);
    sample_manager_inst.add_one_monitor(module_monitor_48);
    sample_manager_inst.add_one_monitor(module_monitor_49);
    sample_manager_inst.add_one_monitor(module_monitor_50);
    sample_manager_inst.add_one_monitor(module_monitor_51);
    sample_manager_inst.add_one_monitor(module_monitor_52);
    sample_manager_inst.add_one_monitor(module_monitor_53);
    sample_manager_inst.add_one_monitor(module_monitor_54);
    sample_manager_inst.add_one_monitor(module_monitor_55);
    sample_manager_inst.add_one_monitor(module_monitor_56);
    sample_manager_inst.add_one_monitor(module_monitor_57);
    sample_manager_inst.add_one_monitor(module_monitor_58);
    sample_manager_inst.add_one_monitor(module_monitor_59);
    sample_manager_inst.add_one_monitor(module_monitor_60);
    sample_manager_inst.add_one_monitor(module_monitor_61);
    sample_manager_inst.add_one_monitor(module_monitor_62);
    sample_manager_inst.add_one_monitor(module_monitor_63);
    sample_manager_inst.add_one_monitor(module_monitor_64);
    sample_manager_inst.add_one_monitor(module_monitor_65);
    sample_manager_inst.add_one_monitor(module_monitor_66);
    sample_manager_inst.add_one_monitor(module_monitor_67);
    sample_manager_inst.add_one_monitor(module_monitor_68);
    sample_manager_inst.add_one_monitor(module_monitor_69);
    sample_manager_inst.add_one_monitor(module_monitor_70);
    sample_manager_inst.add_one_monitor(module_monitor_71);
    sample_manager_inst.add_one_monitor(module_monitor_72);
    sample_manager_inst.add_one_monitor(module_monitor_73);
    sample_manager_inst.add_one_monitor(module_monitor_74);
    sample_manager_inst.add_one_monitor(module_monitor_75);
    sample_manager_inst.add_one_monitor(module_monitor_76);
    sample_manager_inst.add_one_monitor(module_monitor_77);
    sample_manager_inst.add_one_monitor(module_monitor_78);
    sample_manager_inst.add_one_monitor(module_monitor_79);
    sample_manager_inst.add_one_monitor(module_monitor_80);
    sample_manager_inst.add_one_monitor(module_monitor_81);
    sample_manager_inst.add_one_monitor(module_monitor_82);
    sample_manager_inst.add_one_monitor(module_monitor_83);
    sample_manager_inst.add_one_monitor(module_monitor_84);
    sample_manager_inst.add_one_monitor(module_monitor_85);
    sample_manager_inst.add_one_monitor(module_monitor_86);
    sample_manager_inst.add_one_monitor(module_monitor_87);
    sample_manager_inst.add_one_monitor(module_monitor_88);
    sample_manager_inst.add_one_monitor(module_monitor_89);
    sample_manager_inst.add_one_monitor(module_monitor_90);
    sample_manager_inst.add_one_monitor(module_monitor_91);
    sample_manager_inst.add_one_monitor(module_monitor_92);
    sample_manager_inst.add_one_monitor(module_monitor_93);
    sample_manager_inst.add_one_monitor(module_monitor_94);
    sample_manager_inst.add_one_monitor(module_monitor_95);
    sample_manager_inst.add_one_monitor(module_monitor_96);
    sample_manager_inst.add_one_monitor(module_monitor_97);
    sample_manager_inst.add_one_monitor(module_monitor_98);
    sample_manager_inst.add_one_monitor(module_monitor_99);
    sample_manager_inst.add_one_monitor(module_monitor_100);
    sample_manager_inst.add_one_monitor(module_monitor_101);
    sample_manager_inst.add_one_monitor(module_monitor_102);
    sample_manager_inst.add_one_monitor(module_monitor_103);
    sample_manager_inst.add_one_monitor(module_monitor_104);
    sample_manager_inst.add_one_monitor(module_monitor_105);
    sample_manager_inst.add_one_monitor(module_monitor_106);
    sample_manager_inst.add_one_monitor(module_monitor_107);
    sample_manager_inst.add_one_monitor(module_monitor_108);
    sample_manager_inst.add_one_monitor(module_monitor_109);
    sample_manager_inst.add_one_monitor(module_monitor_110);
    sample_manager_inst.add_one_monitor(module_monitor_111);
    sample_manager_inst.add_one_monitor(module_monitor_112);
    sample_manager_inst.add_one_monitor(module_monitor_113);
    sample_manager_inst.add_one_monitor(module_monitor_114);
    sample_manager_inst.add_one_monitor(module_monitor_115);
    sample_manager_inst.add_one_monitor(module_monitor_116);
    sample_manager_inst.add_one_monitor(module_monitor_117);
    sample_manager_inst.add_one_monitor(module_monitor_118);
    sample_manager_inst.add_one_monitor(module_monitor_119);
    sample_manager_inst.add_one_monitor(module_monitor_120);
    sample_manager_inst.add_one_monitor(module_monitor_121);
    sample_manager_inst.add_one_monitor(module_monitor_122);
    sample_manager_inst.add_one_monitor(module_monitor_123);
    sample_manager_inst.add_one_monitor(module_monitor_124);
    sample_manager_inst.add_one_monitor(module_monitor_125);
    sample_manager_inst.add_one_monitor(module_monitor_126);
    sample_manager_inst.add_one_monitor(module_monitor_127);
    sample_manager_inst.add_one_monitor(module_monitor_128);
    sample_manager_inst.add_one_monitor(module_monitor_129);
    sample_manager_inst.add_one_monitor(module_monitor_130);
    sample_manager_inst.add_one_monitor(module_monitor_131);
    sample_manager_inst.add_one_monitor(module_monitor_132);
    sample_manager_inst.add_one_monitor(module_monitor_133);
    sample_manager_inst.add_one_monitor(module_monitor_134);
    sample_manager_inst.add_one_monitor(module_monitor_135);
    sample_manager_inst.add_one_monitor(module_monitor_136);
    sample_manager_inst.add_one_monitor(module_monitor_137);
    sample_manager_inst.add_one_monitor(module_monitor_138);
    sample_manager_inst.add_one_monitor(module_monitor_139);
    sample_manager_inst.add_one_monitor(module_monitor_140);
    sample_manager_inst.add_one_monitor(module_monitor_141);
    sample_manager_inst.add_one_monitor(module_monitor_142);
    sample_manager_inst.add_one_monitor(module_monitor_143);
    sample_manager_inst.add_one_monitor(module_monitor_144);
    sample_manager_inst.add_one_monitor(module_monitor_145);
    sample_manager_inst.add_one_monitor(module_monitor_146);
    sample_manager_inst.add_one_monitor(module_monitor_147);
    sample_manager_inst.add_one_monitor(module_monitor_148);
    sample_manager_inst.add_one_monitor(module_monitor_149);
    sample_manager_inst.add_one_monitor(module_monitor_150);
    sample_manager_inst.add_one_monitor(module_monitor_151);
    sample_manager_inst.add_one_monitor(module_monitor_152);
    sample_manager_inst.add_one_monitor(module_monitor_153);
    sample_manager_inst.add_one_monitor(module_monitor_154);
    sample_manager_inst.add_one_monitor(module_monitor_155);
    sample_manager_inst.add_one_monitor(module_monitor_156);
    sample_manager_inst.add_one_monitor(module_monitor_157);
    sample_manager_inst.add_one_monitor(module_monitor_158);
    sample_manager_inst.add_one_monitor(module_monitor_159);
    sample_manager_inst.add_one_monitor(module_monitor_160);
    sample_manager_inst.add_one_monitor(module_monitor_161);
    sample_manager_inst.add_one_monitor(module_monitor_162);
    sample_manager_inst.add_one_monitor(module_monitor_163);
    sample_manager_inst.add_one_monitor(module_monitor_164);
    sample_manager_inst.add_one_monitor(module_monitor_165);
    sample_manager_inst.add_one_monitor(module_monitor_166);
    sample_manager_inst.add_one_monitor(module_monitor_167);
    sample_manager_inst.add_one_monitor(module_monitor_168);
    sample_manager_inst.add_one_monitor(module_monitor_169);
    sample_manager_inst.add_one_monitor(module_monitor_170);
    sample_manager_inst.add_one_monitor(module_monitor_171);
    sample_manager_inst.add_one_monitor(module_monitor_172);
    sample_manager_inst.add_one_monitor(module_monitor_173);
    sample_manager_inst.add_one_monitor(module_monitor_174);
    sample_manager_inst.add_one_monitor(module_monitor_175);
    sample_manager_inst.add_one_monitor(module_monitor_176);
    sample_manager_inst.add_one_monitor(module_monitor_177);
    sample_manager_inst.add_one_monitor(module_monitor_178);
    sample_manager_inst.add_one_monitor(module_monitor_179);
    sample_manager_inst.add_one_monitor(module_monitor_180);
    sample_manager_inst.add_one_monitor(module_monitor_181);
    sample_manager_inst.add_one_monitor(module_monitor_182);
    sample_manager_inst.add_one_monitor(module_monitor_183);
    sample_manager_inst.add_one_monitor(module_monitor_184);
    sample_manager_inst.add_one_monitor(module_monitor_185);
    sample_manager_inst.add_one_monitor(module_monitor_186);
    sample_manager_inst.add_one_monitor(module_monitor_187);
    sample_manager_inst.add_one_monitor(module_monitor_188);
    sample_manager_inst.add_one_monitor(module_monitor_189);
    sample_manager_inst.add_one_monitor(module_monitor_190);
    sample_manager_inst.add_one_monitor(module_monitor_191);
    sample_manager_inst.add_one_monitor(module_monitor_192);
    sample_manager_inst.add_one_monitor(module_monitor_193);
    sample_manager_inst.add_one_monitor(module_monitor_194);
    sample_manager_inst.add_one_monitor(module_monitor_195);
    sample_manager_inst.add_one_monitor(module_monitor_196);
    sample_manager_inst.add_one_monitor(module_monitor_197);
    sample_manager_inst.add_one_monitor(module_monitor_198);
    sample_manager_inst.add_one_monitor(module_monitor_199);
    sample_manager_inst.add_one_monitor(module_monitor_200);
    sample_manager_inst.add_one_monitor(module_monitor_201);
    sample_manager_inst.add_one_monitor(module_monitor_202);
    sample_manager_inst.add_one_monitor(module_monitor_203);
    sample_manager_inst.add_one_monitor(module_monitor_204);
    sample_manager_inst.add_one_monitor(module_monitor_205);
    sample_manager_inst.add_one_monitor(module_monitor_206);
    sample_manager_inst.add_one_monitor(module_monitor_207);
    sample_manager_inst.add_one_monitor(module_monitor_208);
    sample_manager_inst.add_one_monitor(module_monitor_209);
    sample_manager_inst.add_one_monitor(module_monitor_210);
    sample_manager_inst.add_one_monitor(module_monitor_211);
    sample_manager_inst.add_one_monitor(module_monitor_212);
    sample_manager_inst.add_one_monitor(module_monitor_213);
    sample_manager_inst.add_one_monitor(module_monitor_214);
    sample_manager_inst.add_one_monitor(module_monitor_215);
    sample_manager_inst.add_one_monitor(module_monitor_216);
    sample_manager_inst.add_one_monitor(module_monitor_217);
    sample_manager_inst.add_one_monitor(module_monitor_218);
    sample_manager_inst.add_one_monitor(module_monitor_219);
    sample_manager_inst.add_one_monitor(module_monitor_220);
    sample_manager_inst.add_one_monitor(module_monitor_221);
    sample_manager_inst.add_one_monitor(module_monitor_222);
    sample_manager_inst.add_one_monitor(module_monitor_223);
    sample_manager_inst.add_one_monitor(module_monitor_224);
    sample_manager_inst.add_one_monitor(module_monitor_225);
    sample_manager_inst.add_one_monitor(module_monitor_226);
    sample_manager_inst.add_one_monitor(module_monitor_227);
    sample_manager_inst.add_one_monitor(module_monitor_228);
    sample_manager_inst.add_one_monitor(module_monitor_229);
    sample_manager_inst.add_one_monitor(module_monitor_230);
    sample_manager_inst.add_one_monitor(module_monitor_231);
    sample_manager_inst.add_one_monitor(module_monitor_232);
    sample_manager_inst.add_one_monitor(module_monitor_233);
    sample_manager_inst.add_one_monitor(module_monitor_234);
    sample_manager_inst.add_one_monitor(module_monitor_235);
    sample_manager_inst.add_one_monitor(module_monitor_236);
    sample_manager_inst.add_one_monitor(module_monitor_237);
    sample_manager_inst.add_one_monitor(module_monitor_238);
    sample_manager_inst.add_one_monitor(module_monitor_239);
    sample_manager_inst.add_one_monitor(module_monitor_240);
    sample_manager_inst.add_one_monitor(module_monitor_241);
    sample_manager_inst.add_one_monitor(module_monitor_242);
    sample_manager_inst.add_one_monitor(module_monitor_243);
    sample_manager_inst.add_one_monitor(module_monitor_244);
    sample_manager_inst.add_one_monitor(module_monitor_245);
    sample_manager_inst.add_one_monitor(module_monitor_246);
    sample_manager_inst.add_one_monitor(module_monitor_247);
    sample_manager_inst.add_one_monitor(module_monitor_248);
    sample_manager_inst.add_one_monitor(module_monitor_249);
    sample_manager_inst.add_one_monitor(module_monitor_250);
    sample_manager_inst.add_one_monitor(module_monitor_251);
    sample_manager_inst.add_one_monitor(module_monitor_252);
    sample_manager_inst.add_one_monitor(module_monitor_253);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1)
                break;
            else
                @(posedge clock);
        end
    endtask


endmodule
